`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aux0MJ/nM8JobzhkNxIDaHWl2FJzKzwLdyLERcMkfIplr9BfT8NyaoO/SrbScFvxp5rBgQf3XclE
YJPmk2d1og==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bho9XGrhtNvuF03kjgkL8BORp+/XinWPutCRCx13ydWWEhJVH4/XNRrTceZB/mRgrLRK3BG5/wuv
/zG+/IrJ4NIebBYZWcorfmjG3cKvU5DEvBOfLUkUkbyjogfSNlEpk3JnBO3G3wBrFhqlltg6Wk1G
kQDKCy+sMQ+LJFzL5mc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GG+7HajAGNCjExqpuM1Eq4k6N+D/Pm3SnJVxfdkHmYEKY5HZrpT7+F/xzkAkBePC81k6EA1rN0OO
6jcMzNSiGcC3kNjJ7tosk/qMGnx6T8kdpbJ62kJWDcu6EyvQaVHTs8Cu0vKvkN0UWxm2oo/pxOR3
0TFO1AtUtg2I4BWsyFPGackl75LbMv6uXtjaVl6D+NV/mF3/gHqLB3AFMNgdJ6055ghatyT0N5a0
ZgnrNQ3kRvW49OvAkWySOgW+ZZIfzwPVk5a4bB7FP1sl5opQd4C58ph03ImpEGNaxfE2eSY5/Xin
qCiBeshZR/YRUtNuVsox28ZRZGieb1WjIuLTQQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ByVmYSy8KxXzTiYWM17aRPF7gSoAsinaZ3NzGXy5slXqEc7Orq6Yl99m/UitD6EfOpyhz48e9dBt
ljxJq0OYy+BhiEJjbM7LLFYlwL3eTg8h539HeUwbRi+7XVdptu66QstAJkZ/nEANaEbUE7pYUvy9
d+oC7DtotYxHuYCvfHI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P+hPhEh1kOsWErQXnimtHRw6g2RqfRtSOMKbWz/ZtAC+7osPQL2gQVpeaBBxDVOOzP9sN4ByviO8
zo9CvFZfEGgb+E9SlWkh6inAcd2YhNPTm2uJvBHEQuVXC2NDk+Xb9StOtHxHGQsZAJu7R/Czjj+z
xGJiiy++DbteAOmcXSxAOylZ9RkDX1mYvSZ/diExRSq9qlzrj3aikBY9UlK8xragFo7k2D/DEEje
ZMVqeitkbSrwHueC0Y/gv9/mti6SSDMRrWPEVeR6fXczBPc0GD8PglwfCW5Yp44wwwGl3XvShhv+
8Jt9McagtuVSjgHzxg91ZVmgypyzO9onX4hFLw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11344)
`protect data_block
jK8Zb9PuBCEMRPqc2QIlVkIMdK8vttHJoDXuOjMlJEeXh1soVe35jda5eve/jcJ0q7B0GFEKNYTW
vg3KQRfX8piMZdZWfqCZuu14/RTJ+4L24dvr3dyQQY9lwNpCrefFNq3HU8KdaC2YrsBSbmT/FCvo
wHyekIE54rgP0AElg6VQe2ve6fQHSbiFkJfLHNiMrL5jIshevXm2mm8Vb6qS5KlKQgvuMBp6zSmU
4jXKSIwxgkcgff/JNcm4B3PqAKM7xgLODftE7NfavWlpMmCeHZKDkv6bnLX30PHA76X31yjLeG9V
h08AdZk7ODNpeIGZy3L71o8M3r/fXOHIN87iP0nDAcRA8UPHBZbDWK1chBxH0ZbKiSvniQ9njZtv
Xn78NRVRligdzd54p4JUYzqOad2AyKFRfIfKdrFzob6CPi3WgKpS0BTmsPqRLJYONsbvaAClhaF+
HpSTAtqyiNEXfPzN8zIE55imV+pIkNkWKPcNUb+I+hHy/RnilKOTRTkes4f118odOUsehy0oqYHJ
0a+Kn14iYwPth7+Y0lJjLnT5+9rdjGRKXauAX9XWITG/CreTiWLuwS2WG34H+POvzTr+Ofnwvp9f
10x57jIgTQwL6ygT3GWovMq9pW+4LmKaCO9lzgjI51R7zV98EYSYhsBTGINe5JYdgCWnPEG6Ag/m
RwYNrC+IsnYBYzNL/JYJaRuqetXIyyqvfVaOLihjefsUkoCO63e8ob1Z5vj8TyPYWNMo319twZua
aCZfquyZoXne658rGRNljaVaVIQ5ZK5poM5UGGmHFIOyjrYzvjEbnTZD0g7A9VprEYnpASsd1kQ5
3BnP/LO4mrFAlxh5k5R4cPaDd9GGpqYihD7vg9DU/tkwT1k0FR6wTfSvNl4rnJoHjuUUAZcn0G2Y
NAa9LI+JrM2RzXdJItj9z3DGYx2t6w+/Ad2g3FBmJGcQce47r/G9KFUxokfGwqO3L8bAPTOQnDOQ
SLIbXKfmT+08f8YD53Qor8ndBAicVjoJ0CKiq7De9Nsd+jsZDb0QuywLicMAZ/pz40y//VLwZMpU
8EzPTewfV06w/2trIQytECx8oha24Gs5AEDJ8tE5VYEeK3p7Vsl9bnpcICxp04afTDWqXFp4BCCA
YUxKXefgMdxwrHg6SfPIEuFwpQiS5jWmeqsoI5vW1+3sLCDbAH0RZsVTcVH8qmBDBDOfBJseEhz+
Ox9O1LqSSgFLNv8rM0WiU7dMhuUQKxTK08irNfKWe5M4rpjZfRVz48HkKu1uMpN9hWKD8ifl4r0m
DahPr5Ro7kLqMRPrAZHKZea1QAmEscJhIfHpZDMA4Wg6Locfa2VUe4MM82BNziN8Fh+tRhn+akSj
3PwCPpG5uXv2BzoS6HPIIAZrHa3lKR1rWK1pjc4rfn143l3stsYPNMEEt+BNGRAgbfZnRjgf3bd0
IhAgror+MZuEVs+V0RtbLGtIoVqwcDezr1DFoj94KEHLnaRDUWDShYr4OqZAPOzrZsFjIORPm8j+
qp5x1jjyjD7sa1PL9j6upvHgb1cld6jw44DMavwm+TczEICKF8oNXo2GAFwFaVLtdL8656Y8WgcC
YBxgtSyVAP4fz9H8RlLL2JqlmgDsQyflp7tTiQLLzPaA8eH3pYqgy61z1pu64ykshCn+cRAH7r7M
ZAdZcmMk4SWmo9i3a3i3r3JzAypTqV56ofYV+MY9LuBtSXrS+qW01b41xgON701ltmQX+h2D3bhG
0aMS120ACkg/yznkxdSPim0Y59rdnBy2ompBddZClCZxm/VhIDh/Pzp00OCRTFDOCsY9+W+9g9zN
o0r6A6yOFyG8mq8P5EYBwL+peXtsjzgiEx4YWpXCPYIhiBmMyF5nGb+8usnXI904OtLQQyIyoemj
fztOxACGOLUrkhIi4vqV9Av4yDjBBq/1+2jhNcPuK7WQS/QDPfIuTAfkLnKYLAC5LXSB6H44OzNY
0DPxdC60/ovgLZZX8wPhegMpKqaIfJCJS14WJdvl0yQDjmHAUidPgAuwy2vkQCMQTPGZe/9AN1TU
nztRqjd5aMnIrMhBhui35xi5VNuHKRiGkYfBNJHoBHnuL7qSKhnrc/Ep7hPj1XXjx1GIMP8g5NnB
5YE6DhKSfzxcnBsjbyNqvANNIn/1CzETpsPSzjRG0IL0Q5DzS0LuyV0IcmncnFprWC2cRGoQW5O7
GUro4CvZif7nZbVCMiDO2rWbE5fD6UTClbsAYKr3cDioxh1PAzjIjZqw/jvlLtEgWAZbM/J5mq7Z
YjsseaVKOF/96E0TLT5MfhCYhnKVnkgDXnyEvgsseNpEXOL4nUUJyGkKXMp/H19Xh0z8xbBtbZyh
ZrLYw+NVQM6i6j7sZbLxEutxFlsiLfUe74pNW76k+KEsin/WTwB98LkaynFoAiWEFZUAcilfj2ce
hjV5niJrmmJnEWaPGBA5ZZDualekjlAbBREpiZ5L8xJ9GSF8lhB7tRw0exZYbqIp8g0IA99fS3gH
hDMoNi8q2vi90tvCzTPzjH+MWuMq0P+IhRaROpXTM11AKrzkK4YCg06wvA1TLorb3K0ysXlfIo9l
nlLVc371GqG+VJfyQd/RUYHYA7wB+fP7wKQYc4O2qxabbGQ93k9IvWvb8rcDyEiX/R/3h5bZx8O5
WCQt4Wgzbwks5WObzB6fQE58mCtLQRmNOrRMgEQvY+LgBUeXYP4B2L+V3yfFos9WP50/swh1JdBY
sx9PIPTe078OZUxHtzleIg6H/pU2AQdAuaK86X1feBEhNZqogpGM8M6wV382iqEtvoqd3Vl5BW60
bmKCBP5a5uR2ebxMzD2S98SypIPCeN2puznrS9Q9RXvu9erMp/sRovW8Kf1VbpS1YcWtDgGEcVIR
zb++BHhW9X/kP95iyShf6fgOjkv9YoeHJzHMBAO+as1rSsxCfljguR5SOrs0x2/q3l+BVtDESTKH
CxQfcbVBVy1sIqJknnBy+gVmzuJv34P3IQmvy5L+3aaf7PiJs5vLeCNpDX5gNJNnbBqNZu2J9czI
pvao/lHid5cgVqvSwQkMN0ww1vcElPp1sLGG4VnyUz+eAxobvUbxGyK9JOzKVTk9dbhmEXDfdkH9
doQBoFrW76vsm2NjHtc2iocXW9XJ42BCYOTkO4BcALSX+Bpw51Q9ZRvxvPxU9lfu0dnQ90IZIlGm
6BrKD0dLyGnafsmiB+EyQQf+48cP2QUUATp+clLNe74bKUOG4Z1ocEZYxWlBACuXisZQzZsTRkUU
e5RgAD7Pjm/kyIjgOcExrCBn8oogsL5d7iA0tD8onhckybyRbJcAgxt6MbvHtSwaM0o4z09j4eGY
XSVgphpUcSBCT0/vscOnqz84F+Br3Csek/WVXGSkPLTjyNs5imAMDXn6QNg+Ev7PZtcIWgTgKwEb
MxwiaOVi6p1wN68PijgipHnorkGg9wdrbdusKceqxpFK5owH56s3pkgg3WnRXSbmr+v+i+2EVlfL
rbCx1ulfOWdGFx+yOCkFXAnZS0jK9althi+Ec/s5rgCVVHLQvfhsW59ESDLRmogxauvtm3FoIGAJ
6Ve9J/7ELH9onSF2pcmSrilxXww1uWHGaBsspGdHxyhccRCiBoDNY5mG5HSaf8+K+58mU41KtVzV
Eq8w1gfRr+B+3sW5npgvbRVDrVJAU8Y+icoWm2TbBP0igkwIkbKM7iHmHk4QbGwc1oER9oDcoJpl
xY8ogNN0IX1WjBEdwjUNk2ZPFepH9E4CynKZYzVUNMonFZyRvQNVbJiwNOgydIniojTxmDxW5KSC
TFs/qRrRiK/QKgHFhhQmYMJL1e2D5URgBTMJLjxtyYTn+ixOWdml+SLigZuz7zr77B2F25es/r2s
oGNUjoyhUyMh6vyTvRj3id5+SyiDp5uII35+XJahbgAulICRHkBZaMdYW+p7cUGEeao1kQvs3hDY
Vmu1XuRlJzAcB2pTFXP42RpXXceXNbFst3PFq/W5sHWl6qpj0j5DgLpyJ4utAvoO6kwXsY88PXT7
PDuHPtiRpsiR364jItjdqGH2MDLb9tWhgJyTbHWsxAQFBMZxDaR7oIHhzpe3aLo2qZdU3IHHbw9b
fK4ZWNosqcXqWMGrxkLuJVe2wlt5GpnhlcGKAN3IFXaZhGFoxKdZteLSol+Q7g6llJOcXUoqF2Xg
LnOERTFNwe+VHdrwLFZflzTxDp97059tXIcWh1b5Gtg3VbOVQHPO/rLEVHdQCE8wm4cuKe4rnYIH
nwqPnD4kNdsVZTjc7ErMkz9PBr+9d6nDExq5YALWBXKTW28w30sqXKMbW6nnLrFmGiYiddice7Ai
ftoluOPiHWY35gUvFi9PDec8dnnoq5B4Hh8prWMNe0DKkLOXNsCt82XJQwG6Vu7+isQtLU4efw5C
enQuT8iURER/LxW1pg8zii0T2l34iiLTJA5zbIBCu1Z3+aDPTKsGZqj6Xghhxp0hmleP12RfkyRq
iReVVOba1XqxVqpHAVlYBNoEn96bA64IWLH8AUqJehVm2dbsEOOnSyBKk5YqjnFOAV9GfIsMidMv
G3rU5TiIYKA5BWKCW8BIZK5wqElR/P5kjBnozovKicZjYi+wnrNMnQZE+QPnb4mfpQKgLDYo2Guq
92gnK/hLVlFO5YbwmyRMSJJ6/+i0NUqpz04DxadeTTxhWZ2XqbyPxcb0gdb/rgx7NO3m9xQ+qQab
3FEBsVfSctHJsL4XTEgDT1rbAtkj2jt2PXRBhHgZlyO1m9Ngu+jdOvs+0ebWP719YGTP+E0L1w6F
xlTy7Lc7GzRZTfT9DvztWJtcSMu9Yd2bxNdE2/IJz9Iq004HxlKNmm3cLF8/CjKnbxBVxRsmnYgf
IqHhOoU7bRgmKtmmaj4Z28t/UtXPs3IrN6eWJvbdK4tHc7N1L+mgcMHa35d0/Kp/TtJHybAb7jAt
mZ1Sk0byVXgAS2DvCqc1TbhJaaRM390DCmC/PvzqDHhVeFu7YoMlJSp6XfrK1pf2FSL+aro7eRzf
e2n5x0aAKy6TuZd58exMt1xtbZ1StJPrc2rSyo/4MAmC5IXYk6hAMrD/aer6cgsLtZX0b/4GOiNO
zJHxzVnCRiOeCXoYMrGkANVqW2qlFFLqKTfmf5VAogP04VF75LNaW4v6Jfz1nEJDYjJ5csl3K+Qg
nLfmFDxW9n6IA1SjT+WNmvJOramq5zHQZG0wdCEWPsdFWjEJmtH7AOPjkV9osl4v4prLQUzo48j/
NK2WGcI0oZbxPiwnK9QjjnBpERIH/quqWqCh3E8BaiiCr8BPLNVLMNUXFETS69RjXsbKrz/ftiKb
KV4Z//TaMU0r6xC2HC9HRiStMLMQBfwjVuXMutF/XJut77c2x8HuYnVLvkIxLKtcOXyM2+sqh4qo
5B3L9swVT756T1Nm2HKIXzfGz6Ne1wmrC83HI/NzveeJaZhyp9xAMFxLPXHXqgiLbC2Ee8TQST37
0WIevlSh6tX8uTC0t4r8exOSqSPxrfB/OEs9pXEzkaLQCx0aft7GiCIPtBjJcM238iDkM1z68VGK
0UxL9M38S9Tr5HPKYXaqN1Yh7NzcHaMhfVnEjO0zhbOKVRCssi8S33g3bc+ZsQx8oigdu8apxNQl
2yQiiC5tdFbtyryQo64GCM1+Z9n8qDZU6tnRjcGvred57rEsW1E13DyNdp2RTr+XjWGf4EjfnCXE
He4ZCeG4SsIp/q5D0oBBZUdEt/bhlhLeCrD0AgRkXcXENQlj5vL4MpgXWFaSDmSQ33Ry+52wHeV2
md0e/Yh8GN2dW1VyeNty1b1On9vHHULvLc2HgNL8ZfUnDyY7G24XSpB/WR3eLM1IrVgT0RuHwPLA
yqqGBljeSsHOOctuZNsbKsOa8cLTO3ZppVWe6oJDnwUv87pzEMbIgrycWCzvPks2heOojFUpJ1yy
pLzgPmSIQ5WVku5dY3ZW7EYr1z/fvby1tbsasiBRX0N9tpqp8XA1+g/gCBDF9s85k9jNAtU7xkj0
z/xutQlTrqKI8ImEceoCios3iN74JGP9A8yy75lqh2cfkFWgtUY1vKa93q93vfAQEuv5yQFQmhGd
Zwz7lDiGtrdO8iGtPdYlCKaRPBAcC3sGFbVnYbISo+ekMWYh0pnZujnIBYBd+R9l1HNmw3b/kgYY
QHFFc6JCVDjvwtTgnwqSqD6jyB/ylon2IiF9aSWyBO0igNCN3q3lvMY000WNK5TF0eXRxDyTfGx3
opiQLJgiuNzo90La32LycCsu3bxcargLC0DItfKr0UKEK7ywt+3hVvf7lQWiVQfr9wA3n3/e8lAA
nwKszl+MwjE3aY8KZ5avFYRIuTsYTW9GT54RlFwZv0KOwHe62vvx0W+oBWl0ixIM8c9U3wH/GLi+
DuoYyS40Wp1HA3OOkvPQGGa8GadxW77iL2+kcDwAIUZoKcgcg1p4KKLNoX0f4DSsKsV/kiyC9CAb
6KHUMRI7+UYPGD9m4LUOU4BqmP/g9LDtw2USoOvrjY4FvjkXcBuKmcHKFKCUCwx19rv4WkyW/JJv
kuUT2S5jWywxptYzQ8Ml2vOGOUla5jPhSncJFwRAmOqhXM6xf57+PztFEyFVP0ac4pvJbXPiJ2U8
UpNdFntLDOry2jfOtMREjYiGfGCs/vssC3vJrutbZcL/kHpbl4tDaNtixZcmROCvyEhiNAEh3ud8
5rqJSQv5QxKb1lzQJrxaiuuqww2zhGqoJYty8Fj2Yy9kFNZERlqx0B8kI+GyuKbQGJ+Jp/wnE2xQ
Z3yAu1E6qGLI4WYaYxbJGO9J391Zl/mpw5J36yhXHDru2cTIZcjijC0ZdmKb5TLgCoOhPwaiAXZ4
RTVMxgFYENNpzTL9FSxrD6NNL67D5xOyb9K9sQIaB4ed7rePub2AZp9zfQ9aLTw8vK8EDIkvtnAd
5rHJDR+zUpQ8wKU/XDWdtQpJeJBIQf8cH48fIkFf+Q8jND67LRSalOV4qxU9BrbZIBrXbEhIRzCZ
5ulMlmtKcIBnO/fcijvOsDbgTGUUJclO2Pqyx503Yr14L5U0p91pZcKX1l7W0sVubNtLrEjLWZ7m
//VzEnb4TClEXiXqNQEHvd6nEPsYQArKILO8RNV/FNCWxC7EwhcZ0p36jsUmzh5jJiGwnMpzi+bi
c5NmoiP1+ARBCACEI2qAJzPOvIDLBdzqV1hHS6Y4eM9SqUFV9kbK2UPnGGDhceqhnnvmuj4euyFg
0y83jLx0y++2V/gfrB/0MeO99AaHTOkyQllosW66iLt4Z94enhqz2yJ0y1ryv8I8ChOg3TduCdIh
62O/Lj+mNMKaJTidxh50OTxwQOYpJbOYUW3+H/KRTUK1HYfgjbVKOfEM3jW+iRH00lZvCW7daV7K
7NOamOFpNJsheq00kdV8HFoR01vGbCtOZ4Y6z6UonXzJct4YWmHKcw+m46KjIK/vZougmLSGk6pR
iOblOJS7lm07uDmwUbyvGABSx2HQ1SFxBwWLg2wPMKKW0iXEBw3OhglTfBhdTRH7MITiAR/GLcKr
+OM8RYKjPZ7c5Lw1pZNqDF+GDQa3wYqQ+0R7QP1G3853IQxWjZ6gS5a3Lljkq2RvW/vX3mjrTpcw
RjayTDunAJoLBBHE/J3r1dumtDglWD3Bk+S1EPglBHxMNKpp3MLyDYSZRMv2fkOEZPtcF1Afyrif
igiD8NraH5j6gWPBbFUmXKFgVpcVskYsnByRFOy7UWJpHszr7StUd9u+Hg3W7ozvVkJauywJEJ8q
pUI9VSqk15krNApzXBTKcaFL2WmMhqrXlKdZQ+c73wehwgBXaI+Lb7Roizozr07NHW9+PZ/j0NR3
1ycNh/JnR2RvcDalOBjMQlAhXgCllZXDw9IaW5tQkc0F9WTc/sEK5UxEKVmpk1YkMGUDjPBCRSsh
4TuGaw8+27+39+7DC4M9U7fcoHcvKjeRLVKfanvHJS+1GVgiGmJy92gpsYZpmB8jPs5ArI0b5l06
YO83Pwz1teYo1/ehr4Y/T/rHTaRVcAANP4Yxjw27gUBLx3Q7ZAUvYs6Yag9iBXv7SH2iKhnlM8/D
GOSmJjlObRyQpkfw6TmGdBc5rkRxda1qFNXPOdyKZAKiqXQSaTJ0Eoc+JbEdfCfXW8uTj4SLpoPE
3pEk7fAt8e8g+3e2v4mN/IgfvGdjblz/Id8h7EEvRfaiQXcrEGQ6lzcjqXQEbkvb2pDkXBtTmP51
wVN8+tEYapSwAKTEK2/74qQw7HT87W4L6uUTG2Qpb5n/juaZL7Y37WsC2g+WqMzwx6aQIP4OKDiV
LBDiwvgLkE8XPO6mEQ+VXuf7RVnsnLdpao1ZqLd8uN0a0ABXbQbiUiCibuODl3zH0kvRdFKMHMzL
DLyn+OisjL6neQ92C6JBGrCEzYfpe9Qg/LYZSFL7LnfAQ7/I6bL0f7/iZ2eh65QWrNeMiuYZW+xO
bb03oDz+qChk1ovFJrPkUvV4ygsEw9CzoUgZ1yKC1SHFATi1YgxeJLlaPouyNH69+TWqRzGK480j
Zg/iNR+I9yPI5JGgtvL/DiuS6qDD3bMkMRV9rDHBeMR0l6RdFuQg7Mcun6ngZiGOfw44Cp/xpYbu
D8yt2vtwHqBTk+heK/kLQSJZU6xwqsmtmGVwqZ4JFdreCZOPFHrtakJIkNX0O2+k1sEbhaQIjauh
/BOY76A525P4Sg6zgSAKt+mHddF1bS0VZpVPEAfCLqwtg7qBWbsH+wqQkz+6PI2bCa4tRQxWH3kD
EL/240Xkd72gqDZnXpk/vLVMJ8KeYFcDIkXIoBrEkGeACLFhMER21+iquyC+lVG09gfa2cxy9e+u
SqeJ9gnL8fBw+X5gQtXCckM48iyY6ez8UpgkTQuVAUdGgV0mp6hFXfsiZS/29BWJAimguUXUnBQ8
oNJqd3efZpzn+BvwTRvMyaq/5c67stgDAZ12H48guV8v9utRUoE3ByDqoOtSB38dPqE82+4x0hE5
5HD99VVslHbil3rq7wjSl9wecyDQcQJuMjUr9/Ci2xQKPqnzsVLq8JyzVWn3RVJwNCzQO2Hcwi/D
dxhbcnzrKsqqWm9n1CQsCY9+0SD+L2IiARm13ZW0BZyru+oBcP7Q2gSDJkNbGD0e3VEAEk1SA8iv
Pq2Pr8mdJjXVg0Vg1CgDSGziF8RymF9NaKQz3BWr/wAa8Vrt0D3hemy+7EU+eQIOH86Q8GL4+t/6
eeGW2ncnBI5pnk5pXA22IKDxivkYyGXEOEabnzPrSvw5KDRKz9h+a2neuBnMOLQuhooWSEk+I/GX
S8NWM0Avp6tMEL9R9Khx9FBBdLKrrPM0Ga9kC9Wton4S8FMIj/J9Xu8Rw5vLOL5vQhjZdisGXp2M
mHOPwwDNx3lTWzA26kOlXj5iShlBeWlK9nrKO8B+6vJVhD1VwK3Xl+Eqp6lH38I2RDz+yduOWlZ5
na7qN5oVGsNuZQFNtAgHIdMez1Am633kDg2L6adZwCgfSv5OACadOZMjX1/MhBZu+ZGMJeDPd/ih
kybq1nacJiQ7+w4vWNySloYWENhp5Py+Ou/0SA16iSJDHahlnMVBt7RwVHliZhyun7puDy9N66Eg
SIR51CXwET198fsBPxpCHC7xpOr6o8Dmpeu/0Pdd7H2tpYHhAqt61UnDqMNFzJeKvsY/Gmqvq4tr
J4bsbBlFmUow+8ICAO9IY/pcmE3rvTL2OLQ8v///35Vjgo7ijRTOq/LtwHG7540jRlNt7CvCZNV0
mX7K0T4NUJtmr27rf738mgJMRToTzDoNSNy2oDSNFJzEfDKMRvF1irc6Gd2fbqUi3nCFwHKSi+W3
WvYpVmHjMv198+jEyzd1FfX8aIqhCyroHO7R1q3puVnMnidx5Jx5uWAaBR6Mr0kDkpcILElcM33g
m7pgbAoxwCvlEWhbRk/CTuQAZTEaDHBcK7cWQbgXsefidAt488JUxY1Uu6BUe1OiuQlkFVKq+cTb
194EH24VRwy5UJ1zXBz1Zy8ai9jKUaadOKBBoFnnVFGFjJgja/ChxtYZeLnD0vyMeu+6Te/H5vSl
tUWEw1qq+1FfPEKpbFmUJriEAN0WVZCHEWslhuO/MwcWO60uIxLhDKZBelUdJbAIsVNOsVFhFDEb
DB1LtMmnu/s9StTQwSVjQcrBdYxGM829neSoQrZez2vuzXhXqSlx+lAm2+0/wgYOnTxUGV845exQ
riNTLg6GqwUUOM5fMRzbsWPdW5PjukvlabEFOudwA5RaLOVNTuZQJY346LIF1Efug3U1UWoKxCmb
LTt40YDp6rPM+CxVkbjEGja9Q+/ssyWs2W6i8Yxme7/Mpa3pUm0Rf2+G4QWPdOs3Su72WsY52Foh
4BLXhKnMr34Nsp90DiR4ROooRVVojdDIDFBcivam4+V6TMJSPPT24TgYmFdRpCwCgSf8Jr38lOEn
JfpfAiwrvM5ujxR4+hJ1eD9CkizJqxNChMn8FHnDDHFTiUDzfFFbLTOhH+wEQwP1RLt5XrNlmwEI
gWS5bXZ8w7yTPmXsKh9ZGsc6akOf/8Gh2+L/jEzT20/DRvuARNsNr8QQLHNxD/c9B9JPp4Kal7wb
7nUwl8SNjSJoQqev4VQOWQ7OzZyKiACamnW4kkdwbhwyN6yWMIofct3SDqKMMUjZ9IQEIyS9wXoV
TQesYtq/YHMLs6BLZzzIgMWvtSL/Gbphb7z+YczInYBS9jY/M8wipuMz8KNHH+Fj5S7jlZgYIYI1
g3DAtMa4PGxzREz3koHYEqLLuuCPEnArCtSf0GGYsN2knxkMBohX3kUk1G7LwTtjhgz5rHmV8x/G
tzCUqlHGlxP8sIUe69oFM5X+/rAkW+vjdsp1+H7xWnpcqtuM0FgRhYfISUSMgLRsS03c5bx2rEGY
Y6OMwYjHxIRRjunsQ8b1eqPHzowei2di/WXJpiyF5X1gHwtmM48UiXwVZEVPqYmfErxvv3YRzLlB
M1Pwc9abQLAEUwd4o7eRnQ+UZAZcX7kbLI8PLQ/4dbObm/SMqKoIBLlFgxFTMHgjZfLu0hw0Ub7b
04BpG/pNIuXSc4+BZ4ZBladZrR//yVcstI9LFuT094aDVBbq21sq7DiYx7g+covs11JD9zPni7PA
xIuTFuXYVdHbSTqztkkX4l8gvLmuzu6+JDZVw5pXW//HT8lPw7qc+C8K5y5MULMUX9AJL5buyeGx
sI0+3kUXBBBaRTWPt2Ht5uGKrP+SWwvZKpKk4p0VsOs88qIkfCeWf4i3BdohXL9UNtPU0Z0kz8Lc
tX3Yh0Jag7FTPOPzggsh+ZIjwfEV6YB+9CQs+CFalWF0glQ8zkEYRjCIDDEGRxR1EaXhaKwZ7vdC
P2VEdF/DDi2kq5bl/rwBU+kTSmV8HvDC43jcUZqe9WOmc/GcfFQpbESfjwMHWz/lgcnDIkXERR5h
IkyA1CKa8/7Grct5km5qVv8i/aG4VUPrdhDCwJoUuZ+6rEuYZqc9aEKwo9Q1dcv+ev+qRxWjnFPZ
xDAKRJVg8FBnsnBkr06ujEOxXM9FBIEDdgto05y6kQ7+EYij6wrAIs3meGttEdgd8mhWl8sd4ykA
EtdvZVbJuUGc2g3EH4tpmI66AtXz+7yRIqQ3ESEeN/UBl0d0Kr7jh8YUN+UzSJex/sr1UgJUSnL6
U/krw0/PIiXjx6QkkCINAYnSb7P/+4tXuOq+J1s5u6JEZGzD53O/hT7AxGMW+6yvfc6o0qdeAkXF
pSQv0g5bvmE8nAIYWwMhJM8aa7ZKUrCDpxXuba3le+UzQcdhPXJJiD3ZFV0RAsau9IIHrcRB/IBc
5BBnvDDrGSMOEQOwIjYM7vntcoQfQ2fY6nmYb9ufpwrjBhVLWp8I/Vmrh3g041eV5uMw28351gEC
zndP8kdJx9TF2xRujUfOydCuTVde5VqqQXO0zzBkbZN/X5ch25P+KURj8xSEYhde6nIL8YOfi9NU
x4XZnmjfuejW5UjwkEPsLBtTO2eLoM6wfTCZi+Enkr9PkO+e9ISqrRgoKnCcWOEy9BmHBCMYvg2A
9hV10WIB4orVw5Oz4zscCJumqG5hxDESpNbQVmws/a6lmZ734gZzPOhAP2xnHY4F9O8wTImC3CC/
61FuKElGl4BH/waCsuqTgCFlkZhZSxjKtBOcAr1CPCUNEVO83Di87EEoNVoD9rizJcJAX8eYvkvI
FMBs613/o7Wsgd0UhZ+SaXLKlVZKfpZBSGVqfFjDd/6dCSa0NKcxGE2mpFTrBSjmXuXflejNDljQ
b4zuwfQvMzNzJcFiNT53/bhvs/7pGByYuGM4ZfF09jwLraVnAdrCr1xChgJNK2LsnYSmpeAmfDMH
m77qLEa3aGIjdQHM/2KXYC5spv1V8yh6il08skVC7DOBMKsqc2ozJsX2yK8otdeiYV/3J0sPEWh1
e6ihcPyKe1fWSqc53Z/JfvEgSyQtyaW0v7WDukbzBkPW+xlPT8Gf0+zFZ7ve5CIRN4RkJ1hbVBca
a5l61Ohu93SYYhrWLc53jTPcxaqFDIJYz7eYh8TO5bkDC7TcOVFnQ5TnIsVmCDVEnwuH+CFChC4I
ZUvkUaayJjyyl5FVIbJl8rG8rvdN/kvglqRS4Gx1MVH6Q0qMMqYZRhoIMPBS67ugW1ugbrWUVnKg
/oufGy74/WWFMJIkQxWc45agsRGiGCg19JJJhPWxseTZYiZbuvxaf0BlE1jC6iz/YYAKx/fMAr0X
v4zaHVj1UWwOzrEtbqvr1g1+Um0/oz+PVkBiCfAqkuAsaOnCwZesznqGSLIc5E+xOy+3PU051zTs
Wx/Fkq715h1GOyepZUXs+RhcYlhW/yJgeEUnLobfEAA3V/yOY7YJycjTA/Xq9ltAyKhjWUPFMj7z
AeSrSiGeVgrEeD7eygZ8rn29quzmacybno7U3bw3vnKIsg24SEz+3VshlzjddqIf0kJ7lS6h4WLv
+DKCqbQhyV9qToBZS7SCpigNm71MXdTIomI/oWEBN35gNmmi2BR5rdPDHtFqo/7QYQsCvWXcokyQ
t8KVNSHCMI+csAG1S/f3W8XOKiS62PjubUdrSwwpK08twusVmNW1w2Ze/zRESSoggh6bwjc1Sp97
wZGLCpAe/WmAG9SWqZ2fCJaM2nzvJ/nr4bosO+95A3ozBm+fe/bPJBh+P0HolKLYv1zbKMcSscrc
Yxcquo0YMfLMkWe6whMzhbmNOQopDmREusYPi8yCtlAkT+jfyRUx+Km82S0UsTj++HtnKSl6pl6t
p71Errn93wQijW4sARGFXwkV7rDOoaEKWMLDO0AJ+6urFjl7cm04S8YQAMinUZNnw+9OxJIxLdAK
xie2cY8RaETWCI8ZjB1KiS0bTsUFlCKeYxOgCnYk79rvyPw99gTLwuKbMl5Yyz8ttNWGwz0aQnJA
7aEVdtJ7Iw/idcMt9Gl116Vdmbc0lbhoKMHZw7R918GQBYG11EH5keDPF61YRPRRoapi2rJn4bMa
wxhi+QzfTyXC/U2us2ys09iLd/opdaIgkAmysxMRltwEoQGcHGsQaEnaQMD4srLCO4GLmF++hxC0
myD74g1VF6UCcTzY6xO5MjsxOM3LAFHORuJt6FKmy13WjExSkV+ngZaCTa8UMDlohs88AhB892+Y
RJC/fTdk/uRieetoXACxe3ClqZEvRAv9yXFiNzm1iF84YazJyjtQM+c735lDpxBqtogxqiAVwbb3
B7NzClfbYzKRZlCcnOiGKuTfHKkF+6YoPtbZyExFbynBCIBaK2K2nD2gnmnq68/LVbg4G49bzR2X
f1dNchtGJkxTaHpGtI7j6TUDeA077w2rggw+0uTgBT3pTiSGNZXkFaCqukLdRH7K8n/bgNrCXY6E
gmrksslN+AULD8y0ILeO4HeWCL+oYJtErqwgIOrTOLirjpWqhjEw2Gf84AdZMlwVPreg+J2BLbFD
13poAZbzzbxNmPP2hVKHan7zHwN7bN6X6403q0lkyx5Km/yKiHctEuG6JsHtMMUoGY0zUEDvQuKY
m+bEu6fnaL4dlZGIuI5/ubz5tBk8nkHqveirZrtsfb4LMOfIMar63i/RSTksb1+RE5lspq+UfCnG
gpyPmDMHa+hEZHSjnpfWNhVV/BDrGKWjE0hBBw6Dt377oAan2DhKMLtx7ONggwu02ERlI8mo1D+r
EYyBrbV22iPALgf1LVjtxCW3uf/cQYGI+8hDKvqilvLvuvueAx7HDpY6fbhxkYvqtHiYfB04aDFM
ZpuPKJiYZSkyq6or/vz2S9dc2EYdeb4wo6beRDsdtv37lnHD726LpD0nwpczVBDgin2O61uQ5gxD
k28z8jx3xvXYCwBZZrahC36Ten31WWO25HNCcsCQ30sg13to88oUjZrfwo2Khk8eOTW0hBFoj7Fd
JtJJefQdBiglo95wpkqo5HuC1EFPft/LmKr8EhTNIjuKM/YMvWjOKXnF0wZqVt6ECo9IJWXJjqLa
THSkSmqPUIR2nGhKsiPd+C+6i1yL4s9IbMYoRhw42H8b2Vh7Kwu0xJyyC1villB0RKP0HRiKq9J9
HLituNE5ROT4Y5wlVuhvS8etuifP+jveMLPA3vu7X5U+AFYpHKNujIf4C1R3T4W7jjhSdAe4IbPR
R09vOLmmYp4qaSBbtIBUJGHhGQQgvsZr/HWFP7YMd3FcxxqyJQkd2xNH7Novt+ybUOJMR5ZA9n6W
lKXhujX74aHPgUZpD881BdS0mqYbK5afEzMAZG63Kv/KX62PNFEM/z0XrMuEPLnurNPJGoZ6ugR6
mGGHlhEN7MLUsTK1Ol3ZWxDbzKftMLJY4C0yNENpy7vclR6kd8gp00JTJF7j6OKfalFdHjta93Sl
FcFFGWqn6FilXfkNxpBoBxAh9gs5dudpMg9gWv5k8bKgIhkS/MbHO9LFX4Niia+9qVA014Um8IbE
8sDg+i+NzMMk7b+4wN+5XT/V8cA3JYJuOJvABUhRMq91hX4DandlVbcwj6xH5fjahEaUZE8DsOaP
MJdOSnydQGBio7aYLpl7vhYDi/LyW26/MwXCoPDwRV56B9mfcbzH5ArKl4qHbf+30w7RyGO/spta
+4bLaslHz+N1shWDQYy1Rtm8ZjzA/W5rZMNzTynPp91W9rxN8+rC1ts9D1ckvvrAKaE/G8iL1QvY
dQ==
`protect end_protected
