`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GRrveDVNJiA9foqQYPG4SRHe1EJTYjUZvb/TpWMweYPtxQYL8ktT8+GkgLJ+3BdgVczph3It70Ta
XHfqJipBdw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RI3gNEycAnp+w4sqsFo4GcvyLVybJH1qH0pvPcOyYESXuhq9b6JyCgngTvr8EtFS3akVaF/ghRdu
y26RAylpB8iNRsctcc+dZeZd8xxkJv4KkBkxVnCWkGG6wuAr8usD0GWxbibYsylM6mm5KAXTC+nJ
8huUVeFUfeZdNwfDKp0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iDQZq97kzGp74ofR5502u86b4+ebUSaIXMKppHdOvb09Y2qcFtptGeZnvMrV9xcAkzvgJKB8QQfu
PsSPjL6Z016B61lG/qLidZ8ZfsOPhK5bOzBwkZtCTQyUMk05bKE/urVadLRlWZQEPwp9ipC5sCmN
UKeEjBBeMGDuLERt5RLzruC+Kz7IQc0m/09NS0VwTkyAYh3LHGbQgdHNR3uGPo2QGU8+OUeExZXs
D61I1S2Ukx1djs/zqwKwmeyMjyvtb5t1lA4dRVj2tSC11K04wlUYfMGQXo9mObwP9FlYUayO+6A2
oxkBKi4VfXHd3rsTxsWzpAElAhie0xroG/9aUA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1Q6Ufg1kz9WzNEj9WGyOR4jBmrgfGSbj1AOxfagyWr+Rn6AzkxxvRMukL/9hYeLn9lyomiReDZMk
42w9jqUAivdYNFPSQ/ZPF5lw1QgkIn9eofowikdcdvfZrY/XCHtZen/TyX6YPSbrll0+l+PUqiER
pGxF++cXqH6DXUUr76Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CF4JfgjSh3qgoY1B8rAkyNxSVz0hmvtWNUSj2KqsYj44EKav0efd4fHWw5X2egorwn9oHG7TVKUy
qHX7wokMxQH+s02rgI+W0VE4u9mDgVHL15Qvb3D56gUmaHwqa1NCqyMj7JkqO8upHQr23XyFt2bZ
vGxZMRAO6q++GD3BIFJ+9kc2UBSiCYjNsdiZ8NHcVSiU1ihHIqkgpHkW/JqAcATIwhqHJWJfjtMd
Sc4Jbl6WnOO8Xy9Yxyvg3SRAMtA51G6QmIN8egaaYayGvfK8qm9IH8cwBjqkvJVIz7pcBYaEh22F
ejyrsQSFnMqYc1LgyFgiUSAsECrgu54hj+dFAw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36096)
`protect data_block
x6fhQVwKEsUwc6ZSRsR/GsXUbUsk9oRqggdr/3vEtvFSMWresmXn+xmQNc5oUMHURB38JcWWtVs7
GXItgncZbHWUdn+IH+nMaKl2b/0KsKuFfyLl3dkmWFoWjz66UJ+P36umDF4EnZ1dhfBs64pqGjvH
JnUUm7lk3Z7AA4a7aEBwo/efwBa11rBKDOk3Zx0vb7g3aTPt1hgUOJ0PNaG+FCUpPQEMxb7MNSBB
pqPA7rq7+hurvT2P5J54F8vqP2jD6Fi4+6m+eK1sZALEDfSk1sxYk0VGZGk7b846Wli0TETAfyVM
KSle9bfWqCEHnF+QASnCMSFpT51jOo/o/bD6uJRtj2L0S0wpEv2gU/uQDru2+fvghMl4zwYidOEB
YT4jQgpdixpCUQCbWBgOda0nLWbDneQev4RZr2UH03MDAbaR0gLmozs00n716tji3XgRzon2YbYc
yhh3/ccPCb8qnGmEhI8azoVMAuysO//cjkEGI9ekvRhDzgvN2Lmd2plM6MmfVtzpPxcpbkAdBK/P
puh58YgM4WwB1jcgOJnpfQeeiLMIysJHT8jqKvMGJba5giDnWFjd0YbnW2rPkgqLopUkmT0taB9N
CkaUSR5VgIVI7sOr2kE32rO3bgEjqs/8MxNXCCEa7VteZ4uKfKKnzg4K1TsYCPSxLgoHUwrgmi9+
MoTbkBOyWwdM0XV3qkVi+AKPktiuEGV8DDUnKQwRTXx/6+qCOLaolWFUKph9Rs8OxkwfT38og7tw
VZJyXLogH62K/iGoY9jfjZKXgTGRhQgiQVOOBtYL5kHxKVN6QiT5mq72jMHXNmwqxiRmRaORNfSq
m36V+Zv7Hvfq/tJquAAuImCfwnJzs/Z+5jyxVQ5R86cqZNOQwPgGcOiwxmrI2pvi1tp4MHh+gAJ0
1ouFNKGCVrECer/r/Sn9qUyZSH9evTTNMTSOoZm/iaG4bAc8kaUhfTxI07XHlRHpxseS4O8E6Df8
9+1XbalbTfGmyGWJlgsVy96+MGjvBS4cXZOYmdrZKONtMNhUfm9eTeoFGbWcR+lP3DXag6/6E2DR
gQa2Q2lnCgTSkpcbRI2KihgvZlC45Za39s/CjgsHR1kZgSusxsRSXXNOsEkyqQ3f8RdexP085oML
LiZm7Y6wpJkbbMrfyXCtWVyPFS5hfJemzLbtLfFUROIRmR+Yx8Osy+jHNYRmbuyA4dWwBMSAQeKd
gFdhy5aN5iLR76nhSoZ1kItX3mpkQqBpRlT1WUi53f0iI+wSTPdXrX+w7jT+izr0tXb9EKteHnX5
dGQeNt39k71fFuhChdFV7yYpq87GwqXwesRKo0w97CGTOxizlpaxyS5Jr/V3MpA5kPDmo3cEMlXq
OM7FvzIc2HjBK1OPUQYsc1bB5A86jgDVwtubZy8Ch2wt+mQmBskikNPv6x0tkhtY682Fn7Pdxo6n
k2D/0/vH4FB/fvj+l6+vS3nEhpWEsmqyTmrRYfZlGvbfyU9At4+Jt7h7Uf9xT02Eyf7A9lrmECJN
JKTgn2EwLf5JkvYXUztYmXs+11hWEd/5r10FJCUvTufFF2RPcRSxOMqWh/9oNmlq85sqxNkOIQiN
MiccOlRzId8CpICQw7gAsYZ8+1rPh7grVlfNAtU45KGr9uUzd278+/XttkIu0QYXN8b2QdRoeYsp
p9KvgkpZJbAxfzIaUEzs9ApLhlY5XOwan6GH9JYZ/nyZfjgDYrj/FC3l7xS8eEPXZnWQj6uMgaw8
CX8U31B1z2e3UHhGrnOsA9rb0m20VF3FMr2pL2wUObET/1Bu7CCODIMeVIFbUv+C68IhQEv1YB1D
yeY2XXBu2UkIwOAzdV3XIwMGYrwPurKuzOSPoez/2GqDIRrga98gfbOitKmHHgswIl4Fouqa9xRl
phW8KVOR7ogrOsZT07GxLvShGTWKIJZUX9Wj/jPSZmNLVek1FW7TN0BrhR4YXbunT09bOj0v9Moz
B4KhvegeoFeMi/ka0/ikK2G0zz89IN0YVf2V/eKAgXCUinhaypeak1g5ufiKc2S4NylxvM/2Wrl6
wUndE0eqqtrZwgLH2TSZApHMWHj1LHtEpdCMKhuE+ozA5qqShnKlhFavB4/d5s02W+L5IItKeGVQ
jldUDE1RyAU+AznJ5/+4rfXUbVE02HxVCgtwun/1IJl4udERguTd30rXpnM7f3FWrCuNIH1w9qoy
F9kW3WLF1uS0IZgwN+k4cajHfZT5kZxewUa8mBF6dsKFm2Td+E57HXOkvjoHqv+SVSQEMw5YpAgs
1u766wSjWuOPAiDdGJKvmFaTV0i60eRIA/HLw/tVJIgpe7reyFA6XqUlKO0jIpUH7zN1NBIYIojQ
Ndyg9+NqflTFQgI8NETXa057HNhx3SZ0AkMGuoDfhMLicWX8FZ6IgJDwAjjquAbl4oIChWCMADBS
OdqnjRIvsGapWNvTAGWZNqvEv6oCgAQuS8WUU4IrKJu672NSZ1WEMc2sbioMUUzfWbatveG/U7ET
4YLyChQRpLjhK/bWIM1fMeEHZpC+RTk7eIl1Sz6L8wP9LlYZf3AqdPMqxDMfh0GkAiRmOwOzZWeL
LHMJdbsAb/p0QZSdlOLoScU4cvoKGD8NrRx8rd9KL+GWNeKDo/K3/onMmqjDROW73Dy5YHG2hivP
JEXJxoxAz9FdO0uX+ta5irRp7WhlXpwJjGbtAdYCbZ6RGSWO8aiOzxPI69dlBROkoxXXU9AIixu5
3GELkwJbN5FUQMsulTmdb+zU2v4/vvrF75DTTi+rR21sBoyW0zFmjteB01BgCBU+Tdq4CuEYzEnX
e1RgGa7BoXi/6fJBxttHp3/15YL/rseSq7DQEpBcQ2WKGv17S36Dt3tPfQTGxdatP2E6M5/YlsGT
0ONhhxm/rB0HvIONP5OP74iQzLPy5F5h3+6Z9NRukS4rcalxrgr5K5VdEFLxFvFhZ9dwfcFU9us4
3mIHF93Bez+kJQhK1RuYB3zZiMcLbPIuLuTfWf/NyeSUKaa/DhX9bRR3pJnQNaC+iiPPPZyz6WA0
C+hE1IEtbuDUE537Ret8AWFWX5giNQvKRB0YsACNSaiAwb0PBMwDxFaR0+M7J/QW1jPUdhWMKxlU
BIqj3sA3dV7S9FGsglQXTO0aM9z5XgC9g5LWlAiGQzMbZiICoRyzbkTW3zDhpzc0MQwH5C6UZqcj
3USUJKOZx0lkDYO7i80ZdEn3vXfLFhVDZ3QL2z4UABwl6U9bv5oUmT3U964nr6Qzh8bY2let17Qd
h/Xxx3YPN2qV66Bm86J1FOj1Uhw5WgIl8gqLSmx5pUuJVWuX+9dQanjZv3sTQpxYCGUMKUAGh+w7
pS6lQhwnqfnYOFQv5VWMArB7JWpQHwm8BFvOVTAjlHOmqDsP5PJYNbCzHJx1vgksy7Amyr0c2zRh
DbsC6R5Tuz2GIFPKbzN4uSx0hWLROOm0ZBsCHWgkWeVTAMrlDa1ycUXpX6TBSGN/3XusAuRFzomS
rCjQ4WJux7HtsgpE3EpqHyVYf8LjDiCss/gActga357puwUEOyiDnZ0pyAOiWiCjBgVPKeod78cw
yoeE5EtRwozD9yA66seb3Pj47zCq243krb54lSAFA7Jqwi40UhdrbX9ILbcIN6Izxafbs/q06sHe
SLltNKMj/JNUUxv6gZxZhlR3lrRH0MaTGaK30Oe7xC6PEhof3k965GzM8r/Is2H5pP9FDbPmvHBG
37Y9Bty1MThDRSzT1+EyFKUY017K0XmKQB23YULlP8gFUscMIKJv+KIzUpNHFXoUt3zskTL0UHEA
JXE3l4M1u/rcvrrtREWYJylE6pYzz7vAET9+5eynP2Yb0gumx8tSzffWC0H01Sm+4TITpRomRDLd
+h/H7bBkeq5msCiH5qqCIneIw6mPGVpKw52Bg7yHLO1qoa4CcB130OTe/LEsQrq88CWpEz/JLLfi
AWPn+d+6hmpB6qUJmbtgEmlOJ0FQW9mCWIXAu5TUrp4Wyghg/za0+iLfSOlfIcmEiWhd+sdt66VX
S6FFj+rEM6ziBYMgnsFLpg9dgn+dTSRzgSEXnDeMLmfW6wGkxaDZfES1y1nu2Zg+cACfWzdkk9O7
OQgUXV3L6xTDy3rJjzbRVJ/pQRP8rJUkg4NDAcjhhhpiAa29Ki4cVxDcAg9lkjdYyN2S79WBt9bm
E5aq4edb04EK9Csg9oRzP4AFcLdroMnGGDKurmS+pfLnjFtqMzfHyDcCLTJ6NSGnjsw4VdBtu0yi
kxhGAgU+suupaGJoibr8aBf4UXGz4Np2TLCYHPtIYx2xWpLCtYRxTzT+xfjwZmP/xBYjc6nfe374
L/9RO0X8wZpEVP1/Go8uB+Af43lJWpjZs7L5lAwnSMNxPASe3h6aAUdsdMkacV6Eoxqup5s/hCXp
IhxQ/S1rof7frKF3BN9oV4/cO7x99XBVt7oJaeqqr9pBtGZPGYC88ePdboku5HakpB/Bydshdkg3
DvHxgXCjK17qPKoUIYg17ZzwufOVs2RRpTfhGh1ElWxU2FKgn8JeJ4LZm/eJk3k+7YLoFFZGQmjo
zhBZbVjnqSJI/zunEvfpCJenq7MLeNE+w7uZm2RHzMhoi1ngW9GNzP7xpd6CLIV3IXQz1vqbk9TF
aCr426xSdPvXftTInNOxMn8z3ffQV2GM+CDEiAcbVTcx5Y8vrUDf08PNWocH+OhJ4bcV/V34Ps7q
9bxaamP1+6V4UbtcZjVJavWBKdPtQTscI/QpkiGqfYK4p6n6KKXB4StUS9CE1+iRp1NdcvU5bS+K
svGy2CTJuleOSgVPw1k3rGw5YeOBNiHzfrEE3PTmPdCaNQ882SWjPu1T2NNA3yRZQZke4eQrobpd
13E8xwaP13EM4i//nj4z4gOKkLAPbhCKAjFSQP1tKfY7rCoZWXeOxhlpzoIiJwr/iDzTSYuwXqgm
GJxq2MwxZ1YJnoJc5iHkj2tOKZJTLV0sX5IKJqfBH1kElLD8XZDLBGydwkdRGOdDxamckka+WHCS
9o/O/QvBTngd43tnlP2qB0g4kOaI2z8atouvjGXYqQSmd0uZepUYqkMPBF4NcVX52hONfufjJHdI
aoMBQxWqajVMuYX40IE4YJ+ZknzD31vxlv/VT3sr/1Y8Ecj2SGjTx61zMcgl67riQS5fjWMqvcvl
o4pDaZhWI0dTkqsmU7WBmPyl8l3pC0OWLxHaESXs05/1WqqjEiSiI5HqLkw6XgKSulFixkryzi77
tofpjtmv15Jj9utfT6sOaBPXoUaD0OVa1hL3Ey+WdcPLtsT/lM8ZR1h1T6y6DYH8DbzywVgn3+cJ
INqLnNlobu8y6UoRuPwoUDuJpswKBcQBBTHWChs2liyhO4Jh/VwZI0ckyNOqgO7Raidd8ak/RolO
j8HSW0gfmirX/A/6okHM4B+UbaBGKLhM5yJJCH2pr/J0rbPf92DMD+WF7/p8T6ZgUK/L8aLka+ep
lfZcrDvMsIWGnfTMhmgIaGrHj2wqnmMLN4odpOejg5+Y15O7Fcd7lp4cZs2XwSP3UM4RsL39zQmf
0Pn7awecjhrt02A4nwdawdoPUy1WoVTYcPsLw3Oooe1tib9mUWOz5yReiOohEQvIHjYIj/zDvhIc
QItcG9Z6LJD4Rc2OeolbZnqeGNSNUeTEpp7NxjU+f57Krcw6Z3FL98DD4TPvoUuohnqK0uzrtAan
K/Z2Z5S5IpjR1VnZSKpDYrlLS/CvSQZT3YGE5Uc7/Zo4qh2wiJMrO/TBAhbn3ulbWLre4RN4H9Jq
ks4PJa3ooxlvj5KE+xrp7tKbV9nbX+QNf7n6OCp1/RsBqBu9/a6kKrNwISCveZZcmPMhb4RVeuFw
L7o7unMpHHZx4iifb0hC5Imk8ngFYIpKLkSTe790r/to0qRlwhKKh+rVR4E5pfZDHRap1fJmKkHY
YmlxjIhSz3roSMIChaoExjtq9yp88/UsEYjrF1Pin1hlAodFAezpr9p1A0BoUJtN6ChdUtON8M3v
YpB1zzT3EsvusbPvZTk4bBNSulZ+l4F7j9DQYxLeEkiqiQ8iVtscfdnlQJBTbUhHW0GYJoK/i1iX
80AmwKCod/PuQ0Y4JgnRr/AlNihsSeq5UMJPZxMYSp164/2cQAW3sECdPnRr0lq1uRy3Xhpimpqg
pvw3gVM+2v0yh0XUQNMy+623MS8smqhxzdGdo/f6JqQoaHX0kDy6XbFlmta6MAUxabbSTvyX++n7
XqOkc+YL5Da38+dIRt21rjG9mxbrW+BpszzGm/ypK41Eot3bhKTMVj0LiBg9gaSMajgRlLI1RIpG
favyaK2AOKKFMe0Cyd2i7ggUhGMETioriIjKZl2s/YoKPrmq91eLG8LgkLawSpTRBItIfZsU/JNs
IoHzkB4SibiimDFH/uqywlr+uLrKAZmH4kxRYT8EZyuwoHLuMPK/9xfqmDzxvotCttLk7+BFLotu
wZqqRVaGKvQftIgIpuK1W8OEch1vSuwB5mAfxUlYMIibdDpNDbC2PPLOsBS72+LpdSw1iKw9JLez
bLBFC8oJUscUE/EH3/4PR78qLqAN5RFBkuOv3D2ApDUv8BDs4gWuvMoY41y6s/3EpR/8o+AMPz14
3gJOEMLb9flTBpKumX+7iSZpcHCa4QSf5WXQbeSU+SkiXeEvwZqXr3kmcijC7iX7fkUS9tfipn1m
lYn/z7cZC5XDS98Xy+Y1lOxsZjJJPq2aBQVgw/YS3ZSR+VZNjWTotoHfMAN1gh08RhxxBG5UXsOQ
wY0Kze1MvDOHpnqfVic6GshO33FNRJAGDAMXUwof9FNLfnhgxaVUZeSSrwDtYbUdkJGuHnueSWmV
C+1rbjkSGp7imL+sszNXlRNAAY6BTaF6jt/mc125JhSy7sLrtdH7JxtqzJD0HTsiloCHtPzAHHOu
OS7Vo3h/dEWHwRWud98vN5tlmGFMv2d2d+BrYusGse91lO4El4NrrJZOAjfzZM7Ih+Ugwq8ZbWWc
PMFxC/vAHQxy/wl4DxhJiM1VJp0ifJG+cmAuP40fQr9TiCIda+9u2lTlRi8FNXAwiXSV2LglxPZ1
XZBi16NlU/jvIp5FJNQD+Lp5RrXha7JHloR/QElKy1iC9G8zavW6Hp0qTA621lvi/ebTLjpClY+6
R+m0hNN6AzzscXmVzr6T3H9Lv/kYC3VZpDfzZ0rKMwsZXZIKns06tFDjHAuKDGgDVElDfpXXUUZy
LC3mA2ePAoqWaM7tu0kysVQG6Etie+KT8WRb6p411dU9wpto58+c3S80MJqzgnJ56snTY2EFR6Ie
35+yHXza61KY9rUfnkrnMHg8T1cerQSGEgU7PEhxcSGkWoNRvnNo2Ey2Og4MDJSxzt+Ce45kFel9
AnbhAP/eWYhyX5/TneqdHDtKvKGLrQ6Qz5EPI64fWmxvgMfXe5qweKoMB23TWBrQeXuwTDYJ6kEI
MeJW2qxs5uFOt5Ej6R+fplDv1vyarEcHnEAgY+FV/ItizCW4zn6qPfyJCkC6GtXkm5TVHGWBTwLc
gyrZS3sLLcuy9rx19mlcDAt6oJv4wDhweYZBjS9V2kXwlvBr5skJbMcFuoNn6unA6u5BQNsgBBiZ
VrsCI4AuT+XLsN/ZeinP43Pv/rKgEsLICIp0+9sBUELeXrYWvpW/iXkwXQ2BnqwpQqXn5SauKFIZ
cgz7UYV+aUYTRnP7B8WSlAZcJ9hE0CJ28QGaD3Tt98Germ4l8WO7IHNsrM6oxJJkE7e+XoAX+a3A
d/NjSMDsjzyEw9eKNJiPqcpA6yzKAojSkx+4JTrbfZMmTN7qjuGdUyeJ3fUe5xM3kQjGIDzFUkz1
tF6dPmlGtvbhBiC/2y/N0QO0kK+wm8gNIdTgaUYqrlpukM6pCOFKC39yA3iA5eTgJKVQRI0zPqpH
PnDwTVRa9orgtI5biQ/gDfZl7IbPBdzR/7+9izrjeNvh9pvwCPmNE1kNmQ1Q7W6zbAncIGxaozAv
YXZ462MEu/c0Lzv8r/tQ8cu90NAwLhFIrwkYtIgGcqAs+ZdoZJHzf2VLb3R+Ja99HMKNLmhFxerd
4iPXZvTlwfJWcWAtZzpfmXhoTxzBE2k3iTAbrFVKz7eMmI1Z0hbCqlfGF7oF4Eye8acZR+F6O7kY
B5wIn3kKA3fRIDNI035S15/ArrrB1+V827RIxh9Dt6Am2nA4GFOfitLNf6ERWzA5NXUsOblliV+4
3hjgGEarANpuY0VBTLoa3x9fnWjTKsefV0O4FbHkRxXV/hPJDiTmpCE70HoQ5+DWaQc+ZQ5S88GN
O4DarEv5o18GT0g3jykWabGG+N45eUL5/jL6gB5TE51pu1knYDKQ7oCROly1YRRcZiQ+/0rrz02f
YBgILM/mAKD20CXQJmT03gzukUbXCur4f7D6kWifLJUqu33v36ceUWQrxNg78VBVmhdgUJF2p2py
yBZ8mmSvLwVbANhkcQSdBFZOi/ATJMqXsZRLllmfjSQDP4e8DxS5lxpraruws79QB2vR6hCxdqnz
34zWGpGdoltX/4XOz9AVqsSWkyjh9V3Igjvad4OSUEnl5jC1XAXUlbPX8YxMRnOv+pE7qtXpxEMf
PAjdYdWAAlZVK1sq3Ch2ApuLqdRhJwtjWk2dvBPzeZ2fABWQg0NqaX+uyv010s7rHnyoG1xrpMKo
QlHqDYXW+MBXqnyHCs5VePBi1YCNJpY8q/dMHkGaHCnPRgiXYmQ9ZMYfE8V0LYI/DKCl+Pe/CfgZ
4nAL3t+CZbvNEchvma2lkh27GgDP3cNor7xhX1aWMdonHpke1xedizGK0yy5cK1XEe7XTDN4HAWK
bbh69c8HXNbSthXOSNhdLPpf2OPTy+gBS63n1e9cXVLmP45K3/nhy4ecVe4LjovR8GIlhRBtyq0j
+11r8aEHEXhH4WoTikHxEZaMUe92zzlxM1QzBp1mIS7kBKnemfPOxxJpHjDbORR6Euh1pjV4iwcU
LflkcADE3ShpkN73VPxiCzCK45ukvH3dGY8SYvFItjG2bHeIiqJBk1m92LJvVGns7nHpIJ9iJdo7
VELNDzEfqfr9DuESd/fFTqaly9a+DsTB4/wQWk9FXr4/IXkvmn9d/C9ZbB+/4wewMEMq8bxv4tU1
JQUR0E99MjIKkq1vqcx98MDtLXe53IugeQ2/mUWy6JR0I4WOV2Yc7y6YHKkGU1VD3xzQ+Yszx0nq
XX+f+3jmkuHr3c5RoyEB6tDTOwAk9qWovWFpa3l3OkPvUxZN22vJmsB4yMf5Wo7JP7Pz9d8ycrZX
QgqF8yXgNrPIcWBiFfRYdTbNTKq013A2KRYEDS4sybA8VGzbPY/arFSnVtTVZr0wEqNd17un3ENW
n+R4PZH90P5H/AmhjihHaVDiZJe18v5F+o6nni7zSEYBwHJoB0wXZ24Mw8gzMmcUP2gJZab61OG+
R89fD7M8oBqLRzpJdUKvNoBZ/mPmSYLPcl1GgEWvDZZail3LtyooP4pWoGCq9AFW052dQsRi7xCe
YLYkJUDeUVs2LJL1C+hJLu5FGBkxVUMoYC7b6B2dgT5DHtuAArcAwGr6taGDH1qY0UEZRAt6oFa3
eC2nyRLbGyW8J6PDYNqJX6pIYbYP7UfkEHrGXvf/+62pvbbN26aPeYp10L2eTQZOFNuoX+IGY++X
zdlCNOy8//CYyR1qOGgH4+NRMQXsEmCJtxZN6UX6ersyUgJfCLtjXw3omWBCwGzRiS6JVEttSvKP
rlqr6mmAw6A9tYVaU3lixEHrAG94Fxrnlxr8PZ8bI0WXljrR9U70KOmAnTbBQ/Y+Yr2ANjD9AzR0
3QbaZtZOwpWpTJFkD7EyF7NDwPYOjFX5+NEKnH3pWI7qCkAMPeNsKstY2pPYBDY+OflfLrkSBj2j
edXl84PNzB00lUN79UCAmxszbLyvSE5b8XWy9K5dTrZCAZ8qYw2Q2npN7v6oZl5Lz/mms/+YPa06
j7gWXtBMm+jJYvIwobntBUmCwWrhUCKEfnUbOMSxZa8+kl+mscrq2WVeQogmsh2v1eLB032oVtXX
7Tz/UDWKIN97ygGE4cCBzyMOceowo/opBzwa7yor/RNtLAZvDk5h+QNK53mu9HGF3HDLaoq45/sf
yHQOa9GrxucVx+wt2Z7CU31T8xbYEGZZe0Ez7JlaZTfiFbzq2AIxWt8RDx7CN2mVTMW8IXnkgGbQ
nRCEuuF5KBz8csTjNgDdGvR7WB22pSRq+liWGg8VWRFL1dktjM+/bOW9t8M/s1NVadLh8DFsvK/2
EK4lzQsiavbGXMW1bHH22K5HOh/vTcuni84KWz7HLcjOkiasCLLecYcgP/UUI2F/5nc3NsAh5Ydx
Pd6JUtMV7U0PvSR7zuGoqh0tgYowPje3uPwZicNSfrSDDrMgLraamx8lYQtP+Kt/iDJaxgg9MlgX
5h4D+tq940XN5HNFPuAqInzygf88oL7AYtDDoG+9g8Yq/Nced8dEcNRSBw8v8X9FlF3o1i1vYOMF
Tilwv1stbjO1Ko+jKla5JFYwFTrr8nnFoT7fNG4kGgwedPZz/0Qc6KGYYDRSqDpH4soxayTED4gp
Sh8AFCIjLAPkrPBKq17DEDhbtjOE/NfXzSAmeF25qOcxKGjkHLreSbZNeXuk81yCVo9XS6ZMeepV
Yxh40Lhe8i9xJk9osHkd71RMBOkcGQxEjNMVINA0aajmaFdq+X0oEp3+4plp0NzRU2n0CdVM3sAc
/ehEAvtrAulom7l40o9v41O4bU0c6tWhB4hJg0JcnKFQTp60XRnp+3oXqMOizk5HVZvJVb7ZD0Xi
jttpONC7nd6z4MMMdNnUeLgEM09c9jji3F4OWFTmuRtGFHIh8TA88esKx1LQQmaYE7Li20wkNUpB
3GXlGWz9z7Sg3cmt4ldezTsUcYEHTiKbpyTmsD8AACdpIJeIj028PJsclsXlgonT6MBEj1n8Yp58
zEJv7Uto2e88Xod8YGWEY6gX7OHOQne1eyt6lvIe324J0zb6LGxr4kqHXiTO28a2+eQA47mFacZi
KLgZE57Qmqe7Wprvigo2/18AbAX7waznvV1kFXe5PFt+iMpRcJAHw1/GP3CV2x2x6Rd7lvUiXodk
p8hyJ12cg+a7JxUsVWBA92d60aqECvMDDNPh/Kxg2QpWBbsqFWWGb4kfDcFvpy95vFZl+60CLyor
5YYQNHk0OYngFpnVLrr2WY5D++ZHqe0Op4dPzgPNtjvU25PHnk2C4a6UajS4hDo2d5EiARBJZSO4
kMmEE2X0RyoaF6d5e0m8OwNWS+unIWiwVuOyAObyobNUWAdmh213chwOxkgGwwb7i0rLbxPgCAkj
DLoNTyxqRYaphLLg1kS2D4uUDOoR6m+EYL6PbR5lvE2/l8kH3rc9+hoUhCNv8ZA+BNywQ7dH468k
fOIyBaBn2QbDoEAgtm2Zo+AC6xKl0n/Go3gLnQBuWH7NhYOKzEN/EhiRFH8vEBgqnfPnqTI9/SuO
b0tYdtFQWZ/uHVya1Z3OEkYTPwgawPA0uCHVcL6ZeEDM/5AFBDWehC4wjs+/1zdxNrgLqPT8yCjm
kU2qRM87IeVjG14sVGGxE3naFAlaXOgbvCyCKC9hM0ubVueXuqai+BYbmbAHHbq4bgF8PQ8d0I67
6pNC6feXC9SZY9Y4Gcc4rCt09tvG/3RqtZq8LFgRXwo/Hh5MZNC2ZbNbsA9HJGjr7t2CH8r3/3xj
W5ujBcknBFOq3XUVdFj5IeP+26bKQN6t4tqTG7Nd9sQj4BPcjwCly6vSuDRtDIwfY5e9nhaDVqu4
ad14QvmJJs/NSsQ3sA/JXw8txHmITmnu/hg2zr8PyvxGXBabe+axySkORzgFjgjzCa+9PZfkeLC2
jhu8+IJl8C/wt8m2HmhCVymb7C97kgmBjeD+4Dqb9j29qRsHXfZLeImO1XaLboyvIjR/0zg+7+Ys
bPQhLppIcBK3QBC3e0OOYuhGqZ+YFwDZAYdOMYFDn2FNK6UhhZ29J+5NTExZHTDCoaLuiApjmWBY
MuxP+gfMkIIDGiASGaqOTpvr8A5EGY4QakiiTNANw4cZlwwd+1rvsJz9WxnYmGAEXvjGqGfIsjdd
XazXU2I30xvkg3zAIpqAM/CWm/r+luSGbN/4XEY+9ENsMYgmogDb73JtW6pyUmRXE+TTxlhls/Cd
y5zDtw+CLZOEBn2Q0ENRN4bprfhoMmak1bkixUiuK1cBKYAB93KNJaXXxEssvwvQBppAKakggptG
/6/dofzzOvTBAk+bZGlxc8ZpgYAH8ILGVKo3VakC4j/1lHZfk/a/VQ8qfUpQAutdGdfZmWdyI8q9
oO+CXAaaM02NrFw7OTVecuEREUrEwc7q7djCWqacAhYgE7VkqmuRjAnvFP4rp1QP1AkQKaFuAh6M
ihUIOQRLeiGqwBwFyTR8gF2HsZ1XiN+6/fgDYy96VqK6OlleRSBDbzL9M1EQNd9UeIS9HTaxnbQC
pJPkgkfB6VbaSksCLJOMZH4pg69gJ94cye7T5M6Z/u/lH3Wm4TGd7Y13jy3N7JhhSy5Rk2fmg2eZ
vl86eEyO7+gRfFnwyA2B5G0v58I67YprnxqbSovbL/wDiGYJg+0poz/Raub/MfDkvadjsgQGu+Bf
gqleR40FGmhEnTWGbT/RXUbYkjTyu4HL11UL0kfyephVzVKTJFpudPCg227tRVWe4AhXnnIBy8PT
LfDmUYab8h4hEdCxegBsuXX5qFunDATJIGXqFpWUN0hN1Ey8+1prGlAtbfWsh+7XAHke05/G0v3k
poQ3ihm5nkgyqE7ZcFBHQJnXf7OgkyALkwl6e2fIbBMqs3HgB/uaLgeOtiFubadQsm0x69A/rTXL
8hoQusGyiNmt5W+6v8BiSRZOmBHlEE5WlBl8HIl8nUImPZF8I5mhcSiXriQlxUmSSrtGln/ZjRZK
iD39kI85RUPcE2A70NgyzYGH0V8F+YalPFj6IiDWQlPkiwlJRq7ncpV1L8VTvG7clKUTBbhniC6u
V5QjaWxTLwlld4bnhnF6uiqvv001/ekm0nzkUYM+6fM8m2WWgpG9ldNTLxR/ZzwramjFBh2J/e+a
+aEDUApcyxAYxhL6vCbx8EHnNt8q42VZd8kwHbEdyB19/bDOaaRr1f1hPbqOL+g8FZxm0gg5nQ0k
/vcf7SAcCt9acMJkf+3lCtHzfBIP+FJ2g9WMnj+jivbrRpd8EJI7pRKWgDK49N/+uJpCQtSlRRj8
qFUaJ8w/p59ileFbxrXzFW7FdjI+xR59F8E4oYZV+P87li+qDqukJPApOH7AHZeSGRi9p9LNllXR
aJ0LfpLkVzMl6wmfC8JCVvCMQU7+jr6C6Y1NArjradp6CNhQyOlzdGYZ947TnHA7t8hm2VrzuBrq
KpiCg4NNDv2W0142pNsun9laTf/m/yjRHVxn075eRP/vST8IgEz7eHMdtPLRKUoywAL59kutismB
x4a5LBOVib5uDVqXG+OMZWRQhjudGKCu2YcB+zCbO/HlMODRw2kvGYr+EUkdzW4jAsjpPINjlsgJ
2p+rWCsWWBkJJZ42L7tKyyOzMMofK3icZ82KwKWYAvW5gjB1NPfINJAwuavykTyix/4sHkr/NC3j
bAAmeKJHoRXN3wVMdU+ScSJ331nd+qvInzs/z61ZFRGnS7GKvXrl0Dlkm/eEJJjk+v1s5pIZa8ZJ
dG3esJrTEWG0ZsDYIDGc7p15Frj4sBoSKBC+D+jVzhOqqr8iWzPJkv3vXrKYR0PcU42JJ7166pET
EyNJsLw1fhNsI1wu51IGKVPVjlPWIaf05V8sAikozJ5KR8RVZmKgkZO0Rl6V1+j02016yjPRS0ba
WypjW0M9R+eJtyCFBfaVDqH0wShJ1YLQmMf96ZVg/7guqDxy4gMtua+69CGskHwo+xKoZo+uoJ6I
awEspksV9W+SXnTo8T6wOH8Acn993b7A469uzW8zEmUDiAAZPdcQy6qsaxIpY8Vw8C63caPpkOTR
lWTd58HgNomNwKCYbDbf6J9CADzQPO0SMG1AKjwM00mh1pNbsCJ5tSOUs2zUzvLHVkHdS75pqhRp
1tV7SLDbiXO1Vwd9XErExm5jPRFHItmsgYdURViclTsVVSCxf6B35t10nqcOA7CVF9fkoJ5CB2gY
cLrw6fLlzuTV7SSgeTC9M6kLfkIKvqMtii4oR7nU97IQmxrVkDbDTDnBnCQ2fGzQse7wtERJPnRs
Nkk/TfjB5iZR2goX/twsGavBMnb9U+S7gUwb98ZqvIZW8gnHzVdnJ2BgjQq5eL115ddiKoo6oCKb
+PDo4c3tPLhiostKJEQ8F9fe9uLIRCHfz0CJSgdXzuLv7URukHaMkdui7j8boaIfTMjeB2GDpj+g
uZU8Qegz/7t5fwhuXDHGexb9/7ccRtSLjP8IDt0yA45UxyTYQvJmUauE1BLJgNeMLJF9eSQh0loO
4fQV0RlIimcne5m4OKnDawlOOjO9mDXomEVhIBsoWaxjjohzH7fWsCjxUib3AUupIF5Oa7xw9Knt
ErVHtsvk/QeKLyWvoMtEXVGVRCzQqSg2b6wK4rDH1IyFJHsrDD5SdR86ZxJOEFDE7d341qTEKchI
MEhKfnIKTTc6FEnzcb5ryzY/ZPu11t23noadVvBzT/fi8WhfaRMMDdhqkl3NBalCbngcYVjNiHek
kQnHl7z3o2Qowp/DV0H4pxwfRrXxOUCSmuBhSw5+iujB+zuNEg2BDFPIhWJtLlGuabGIB5zMaCD+
ejUmPFF8I/4VVrRedKjIQeMi0idz7YrVjVVN/H7ri9tEA0WsIHdTcLO2i4EvuWEPh/IExivqbsh+
chhcetrxaZ/T2WTcTWHC8W++SlBV1jDkxkiHUkeHAkOG3HQU/pzaW76t36SNdmIUwMxdFzKAbhYm
RzES0MDDVHXQBJqvxaTQ1IUfGf9qsAzqciA9XrsVk2D+c/IIucjteFrV/mt2bz0GYopS3dHEs7AY
o8OlFeqZQTxe17k7l2IHLzKSO5+sy7JiH5WRH+k/7E5o9BFwTGk1+utXGBEM5vVxrqSreNptRkoo
vTkSWN3tmcocI4Y88SVxZEmIYNN7KV1ZhD00zVvem4oBVefE1LFmHMj23opdp1Yh0dz5Vf37RAV4
Uq3QgZWu5DzFLTZQd9Fly9rXPxpkiYYe/iPIMWzbFeWRij7aLMSqPTpu8NkH9FXLZkSDY4703eij
UXtx8mLhJ8K1P+Cf/FF9+6rMmHdJ0pTjbqzkdik9QIDvWw0BJzDRfe1sIvyeN0Do4g/7RKNhs50X
PmWnoDhUysnjFITW/B2H3Hxor/14vOBTDjDZ+fZIRg3EZ+Hh6PHq8NF+SIOm+UZlPBZUg2/cVH5E
5nw44GxX4grOOiXQIfdnom63BQ/HTnANRdjheLWo0qVAu8hM0Prgxc6AHiOCVC2B7LZn/5EPFU7G
Crel3AoPMKiUK3RgUNSQdcbQAsewlMGxGils/DcY9v/k8VqlPKM8frvLkP4/hN6ezdow3nXtSlG2
dTmENDj4cSCIcpmLLhBzqjf2tLj9Z1SjVugaKHQaU7V5xJFNHG2BWfXQ5zMkn32SsgCfJXRBO6Xd
XPKNB1d1lQrb0y6BI2EfPxptZU8QpzZg333ISQfY8Ay3Ko22lv3Oo6C04kD6jcEDBDjjwWPXisMX
spyzrg3vp3OFcz4IiJuiABvSFbdWvVkooBAd1NN2HPmwXRjBsJJuF9jaT2rLsV6pCxEdI9ZVnXPN
AbIj991CTch94vT8/WK2NOmPk8Ve8ajKsZUMz3dUfTtI6HYmppaJx7UUD63bqd07mOvAjRW9rcSN
CflLM+bIoac2g+dH0asphwyhFofa+TgDH3rLwu62dIMZFx9Uyt1BJDprr6wYEu5kim3jrckW06Yi
VEGwgBHVPZYqnL/ETDsulU9Gy+ErKwNZ1lA9IBEl8b/xDbf3lN57er12icPPjDjkwgq70NcuQcI+
qT3Y9F812e2xR7oneOXKU7mX/ejMWY9NVC0GwYjl0Of1AKinv0jhA23kdIu5Qi8P5FcU+O8TEq7U
zKbrLPtYl5EwJOPgowr4nhhos3dm3U/f2xzSAAtIbRd3xb3+JQkK/qfSe34JKFLFpKIHlSzydDVg
rz9mYj2dEu9mLRj4VtuNq0BAwPKzM4P73zQKexsJUz+aLF8EWXKZK0zuKnOJWWdczueCftUOkfOs
maIGXg+MiMzTVb38Mru3XYCaftP8xGAtWOSGFACPpO4vU0ft07iv6iYQntyls5OHyAAQgKqlCSNH
4oU+46WKdph2PQxvxH7sH7S/aTH7otd8adKWNfDlXoLvXBfFo1B2jzhXPCBWv9w22rPJImQp1NEI
MwwpvHCUI+ssuzI9j/BhcD1EwxOG1QdMQtR5WH+/I+j9tqV8QUmlxYcIyEXGLVvUjhQQzkTAxowT
mDGiA1nqO9mdN3NafxUocwPce5HJwSscDbDfgT+0A6RlMOy8CTMIOVUEj4e59/tXoJCYuPEPsjjz
jIwchCxWVC52NadzP5n7ijjkdVW+3j0YwQgG2jwhFxpb5ugVBwP3YclTUShMjyLFCpIs/vD3c2tU
FRhQIn+UXegWsZjZ+oC525oQPG0cplpoxJVMjog30+dBdAZKvCEAoOnUjedI48c+LrQBxtmKUrzK
WtQJsx8QFywnLGz7KXAXZrH6d1QEpusn/sDs5xXy9WXOj8dcp8YvqlV6w8F0coKkm++X71kH9YyL
i0cez3LB+8I0qPaEGBBkf6ask5Ud2c9dwiCZTm8SOAv0IJKhdRAXttxOLuXYTvniZJBMppr9jPgL
pNv0KDDG1vR7NfvCR9Md6F42zdVHbI4dWdgwt49Ua624qcY5GyFkTAuCv+STMnNOCzwhp2An8H9H
tLDO9nwjVbMAaGPqAiVl8hovHKri4FbYZdeJPeEwfzcxd6tYj69d3PCdfH9MZb1tCuyEZ6eGzs6I
Aiag5pbAdZkoo7JUy/Petram6OzL5ev7dqIqCvoRIYvjG1SsgQhzGmqGgx3VX+y0rFRzoCuDfIOK
UQEYHz0mty4YxOZdi2+Azwom2XxmTj3/Io1avPWJOzRoq8ZoZUvKuRtGgWGSxejFp9x7wElVSUbe
yqXTBzx6H5g5MZfwK/YWHcXLMH7Vm8TGBc24iqUjaJcQAe8ctgsBOmAo14/+3ZwIVEstSFF/l8Hf
bII+I2y9EZSgdUrOX4RQOEbtofriFbHiXbS/dLs+4WSM1kTzJ4k5CMNdB3ilgUUko0Muk6sUahKk
ClPoIxiTGXCFk2/yR6+dl2zxjj6T3UZeX5Fr5yfZPObJNfrNuhBxCgEsrCZvGJdcD8gjXMkyve42
RT1xKSf89e4CHeSWDgn82iK1nzP+Cxfvvsb94gM2BwYoHLaQMlcTyDyymIRoeusDjWARiFELSVlC
2PfUeMnVXG3hfrWoIOJcASSgNXAa6zU792RgE+V+cY8AvH/ZHUn2KSsY5/JDucv/0AS+g4+L2tVj
Iktm5XtNDLqFibIDn1vw1y7QIBFXT6wsWhJfysSK/dtqbFqgtEFFFV8sVueGHQ5W7zSPP0C1nau1
aqYzvAI0ZXy2vxNd2P9gN+FNvi1Kd7OvMmVEF9vtdzg6XFxXp2jFgysMYYynOx5yU99srJQ0ciTS
h60Ah8oldrYUdC2OdJyHsjaFl8gvOa+JhZy4D0dj42IpY0OZyGkd53MSdyIIUIOImAS9BtFiZF8T
0bEeB6qh7nclbXfvn71A+VuoFJqoEGsFTouXALyy8kdkf4Z5dX+qC+5busNVCuPhn879T9umI5QG
qZfQUU4ScENb5WfQ8rMwWGrb3Q/k17WexAmqi6WY9BHRQTv5BdWOxxzbGQffiPY1ix/wPbq/lNjt
yHMefdmAl57WRBFWfCB4ttF412165oKH1MBOcxgnXQZfJjJNKAZVjtTRcsZrVIVYYdl/uczqWj91
qPKer3iztUO2cwXG8cWY8DYidD5hs8Yow2kfPqDWljlufqe6z1r7Gtrw8+3DAe19SsAg7JxSZr3u
CEIlwD9F4no02C26kB7AMA58Kaz0qXYZOx6CNaiMp5JOaWk7DIjAS6+7BFQitdQXuu3CODtmdjyz
DGvncNyGmCYUdDZ0MhuX+RU8ygbQBHdVno9KTaqOU2Qg+rOXWIeyBnReWMbXf2M7tfUiRXNPDRLs
PAEv1M2V+ArVoBYPIAWSVTF6S6TSfqQBmDYp+M2oitX2rKNlGxe2XIzoImJX9TI1iK9Kx7XwhPRw
K8x4LiiWH1jEDBUj43BiRapAQVxBbXYyJjb57sG3SRjztrzHOpdJeo+x4hBr/tYEctyH/AaUA4bv
PjwkjXFuGSB5cL5YJnfM7sVuUSProV+LXz/sY9ZOEwGF9gh0CgY9+23nzlygokqQoFOD/PZTWpfA
Qef7BcsHT+7fl/t7Big8E6R0yp1ZJZjMqQonsxWvBn6hvmFLKVW1kIrc5w0kCcQhTIPSAfrlbqqp
u08OGYwGrL4PCF2UhzsELkJAgMCLJS0zq7LOWB3Nyl4Hhco0u7BuMquiPrDQTMQ6BhPUFjw18VPC
f7UvJa6Ph7IMoDH4AnGJLjXjcVh0EOTTlFrDPmigYQg+x+XzVKQRKQbGjyO25U3fMoMjgP+8PPIq
GZcIysyjpwk7VLCPSBmA/j1o6nBcna/mRFI5lFDVac73zqN4p1fY1XjERI3eGKs6NdeFpkICg82f
mbBeF5S9zdcuBQRgWtKe8lI6X0K83pZoGX0NK5cpBmbvK+nkRb/06jiU76KZYY7Id4L7e6NAmfuP
AY1vaSPjQvn742fj0iTgJcGoxxwYQ19e5xZtxMGTlvECmd5eDBGc9VpFc//gjC9FDTElWa+/6TsG
phP/x4rxW559zKaahLfLzmrJjm+CrHg8tH6Op5+nvOIcyhMIk7Rf7bEtdZ6HSkct1ePOhcHcmOQg
ZOy/oS+7a3i9rEQYJCcsJWD3iIdm69HyQ7ZWNWzOqtHafQNzhWzxP3QaJIuFzmWONpYlzlse8YC9
ltEhU5HmIrVtdFdvbou9bvybqmKTscIoGvZQ4BB57QH+3gxjEH1hLXRWaGqbqiNr0BFA+RZD09j7
1lQu7u0goZOKfduz5mz0K4hc7pKBBu1JWJoo8YMVww4Fcqeg5SzRpvyUcp1v9T+yr70RQ6TIcT4W
9JFkwcyI/TuMI57i6PlrRg4DHQi+DyR3gJkg/1yen+s7krxJBgTOa4+wZIDW1JXLAR5LLo/iTTkM
5VgTqBXt+aGHO/N+6uxNnBr/F6wjHmhCtJUjYA3sXkh++8uO3yv6xTgVVG80y8s1FKJc6k4UIUxJ
OZ/VVT0kZd32Kj6P5wspWaDk+PXZ69y1D6PI0BfAMvjie+MBn0AvIJ0rPtRLx5GZcGb+/4IKCiAY
TQo5PI12zM/kq2GYKJo/yExk6qmmzhKz7NY3BbOubEbsfJ715Vvmbwgx90RInGt7u4SHrVgOijeG
oFlZn/lLGTUn4IruBrqMnzd4fhZhBm0kvd2NAqEDtIfQBCVVq2UCdxeISzSlwM1L1aDsV57nArUF
wt9ffbFk33/jWUJF/FzK1ul6h3gDuL7aMo/Z4mDxrqooj2xlLqY/7TDpJej0z+U57bKDoopkWgIS
MOKTRMuwxnR6/GdqqOpIfZgvOkMkZRIfqA4bDAI9+hSLDeblQXftGuzpH4o8BXZwEGwOtEk4aC0L
Tm/ke08ZYHM7TaXyaHxGscHhekvnTzOurQMZnWX83PFilIkxDyj16PbdwAMdyb7R5yorP8muybMq
1Bv74gouslHtIczMdFvrIhJkoWcm7Nzyabut74+YwQgqtLKsfzPrxrHEaoh4Avz6MhWAHaRpDRm5
iQrFfAa0RO2/H9taUWhWhuUR3wEO+W7Q/tFqax1meyctNpiofr8yXQG3RMqvwih0B916n5aCMqCg
9N3bXUAE1J5t0RSdn4SVa1ddLrb6tQOP2xcvBKjIaQFkh7pEZEmZ0fi0pCxObr2RZrJOhYc3Ll3/
dSVjcOQmPkrBYD6ereEEaaFxc4tKVjT9Wats486nozD9NhanfEdr87UaRDnDLmxKMYJJ3QJ1Vzs9
uCdeVteXDOOiDLEG4U2LIMXWoeqKbhtmox2mLorb7WP7bt2uRptLewV3khE0yb8bDVvXKNGmlCnC
2sduc4BSX0jBa0cRpPy0Bl9TWIr9wOg6ADZIR7wZM7lO1bQAxxdQ+UYDDR9bqwROhUBHxr/mLdWu
R2/EXfLoO8aGIMASj/F//SwP+3vGMZWlIFuY0etSDU0+0254ovgnKIUQ/qB4eg6efjZSF6Bw6Z6G
xK+Onla5xr2JhWDG6jnwfC+rQy4ft72FhhBgSOsKF7xcmaOKTDuYg4pMZcHjYAz9vpIPYwXa6JxP
IxRNnfE64aBMYKGAX+CbpigYzXV8QrpX4RWz0xZv6JmaWfjNIJhbwYgSmdNQg5418CKXJ4wWghfu
TeUtXHR71Ie9ClMS5OghCpCEqY0Q5AOxvCNtLkOfXvdNK3Ld6tYtN8BN//Aw0/VIY1ANSL1cvspV
gsEjd5NL3jR2VPhgU1SPnRONEUtupMP3xg0fDK2pKJ0g0XTt6ExJH31NGxpQdysbXPo/jqf49j2j
sb4/NEMxMncgWmM8duYw+peyuHDScP5PWvaYZya+qslIFTUPWBiTNg3oWR+CSO4gevl65F9DPfAX
OfP/h7VyNHFFVV8hO3I5TOrTCRLLlL1LlV3+C1MhdR8msr05zROXRswAcgAF9jXqg4oIHd4Xy9KZ
Rr2zwdsYWWbV2LVheVgAXJcCT5INSFNdbbd99feYZWq5UCDY74fp7lo25qNnvEqXMubHFqLuvDVr
RcCaobFzGdW4wxLc/GlJQviIsduiHCL+MaEkcWnbgZ60s6UST2DkxeEHh0p7sEq150NC5LAMAdOY
NrALb27NvsN/NPpYTRXNaFXgxfvZfjcI2Bzje8APeE06kBdrVPWSwiRR1ZUCDiBfg//nQsyWDLo2
CHHKoRBfm4YEXzdxwvvn0Im5aaB/PK2wDHEmvqWeLd3qLbjIFt9SsyuoJqSyYXORomjkFh46Qref
qqwxR6eWv3U/SCIdnVuQaBs57kPty/Hz1Q6L/udT98l/Yu/JaVknd13mYuLRh1IcCnCVLN8WuGBt
nkUUTlI5OlSsdihx4Z2T3yHnRLGNRDfp1kTbx2rQwtYj6vhxDzYWhBsC+kf2ZqFQazAKMHdjraot
xYYRKM25q9I1BOneRPydktvDHAQm1hOs3j8aYkoAa4JerYGOjI4PTHPps/M+iMJGWtnu3qwOuuui
vTiTZfH3Vqgg8efxGCkfh93a/2Kqi6nttyRauNNCGDhr8327oxAcRJnhyl6PBi0iew178JJ0h/SY
Fiejoaf08OrRPDFZT71xexybuqBkbDoWGuuQbkNcUBFrVKztuJDFT/9K6zTm4OMkG+3Fc6Z9OIRS
QBDq6e/I0u1ebKRanCb6jOUeaZBOeIO4BfFB2TkP76QoQMMoLnp7OHgoXtYTLbZmQaX4IIyKpYIs
vGhUxTx+x1XI93jToSN6YGdGBMl82SQqsab6wEHU/KpnbWlmnNYy/0zU19FB/Ho9MRgl3DaTV7c1
R34Mosb5EaO3qeQi24hk4Y4h9AvQ7AIN93jOR86tp5cO5YryWcDQq5leRz9m+DCgUnzD7/1dgE/R
uKKb2Zhr4p4sA1xs7JG3rVEJ9J9ls9GaGZJzrWnDhj2u8qnWh1QowL87scINaYjUsA1qYroMACDF
Iod8/2r9yNdEFAW2MukMoaJYGVbzOkGBCgN+KlzaVPk4ki9yyIDHujLebpissNFQ4yKt345hildY
byKQ5jEF93uO8VOx3bc8FO8e6a7O7egFdMm3300pFkbT0Q1/EtgKCd67rTVDkw6Yu5MESlUmOfOT
6uXkkkCWts7u5eHQFkGWFC7f9Fc2rKhdqaJOmqxthAkmDi45ziYMEeLxeIwPDJE08pQvcEdIVXma
gQxrIZGDSncw9uSIrsxtlSV/fVsy4obj+HPUn8Ygzb9Uoqd1J72ZaI6o/5BJ6DbxHC9NDU9B2a8R
Kgp67wgAyhG0Ory0INCC0FT8pzDXrKPHtGmo9V2ySmdPHKPrNwgweo+iYeMfS+fs5iwLigK+/5ne
lG1XXJ/9Gl695vj97yzw7i/iEAHVEqgLB/HLv83ZyzDg1iEGwht8wGKh+ZHas4Y+9bI4DXt7D1Zm
gIdJnyOKyEKYJk7u1Grh/mAFjj4R+Ku2PcfCN5jhG7hGqYWh2YjCqtvxWdpUgfp0TS+Fy8NFgQbO
0wrsUDghS2efU1m4NEkNTKxa5wVT7UMIFuR4jkkIMZIBtNewf9nxNyekRQHquCpcYisTVOVb5rCb
Z/KSA5YcFWkH9S8BMMMxVDVyT8fi143sMS7uFIrCdtPhP9MLO7fgd6A2Nj74IA6ROp3VWOp3bAK6
2IP6EbXVdobqyo3SPG56VJaVV9Dp1P6UH53Ueh4ULyHl8Yfe/mJFnUvMetyGE8l0+i8dSI38nEy5
KTqsisPDAU4r/4a/iWWodsVFNkcrezRWOVgsawD6Uux21yMARX0e7h84BiqFK48Caxa0uXmkdFVJ
0KiJumcim6FFNEs4oOfI3e6A6+y0LCC3XvMhwh6oJ+EYCWDAl2PuH0LilHDwHqN1kxZidVcX7HrI
yvKThoOqOyagwAzuRI1Tb6dcxpYLxMADdX8BjmJxWuai11Q1qBXItgbNKShy0Mfz8WsNQAEzTIdH
TP7SxAImTWOREFxCvyuWjjHfEFWe/6gaGTF0tIPSorwjz6Kj9WCU9QffeHtlcmwqgpgGnPQskHoo
lcCa170nQTReXu6MxG4YVsmGy7pmTmHNCF9a92SPUIHZ0ptT0zb6CT2I6qQ//HUckOvVt7x1gtKg
zYhnTtXM5C8kBAsM0fM/3J5UsisJzIfx8IVhuk2unx6DJgC184rcG6m73i66YZaucQNhWafeZ/h8
oVL0JB9z9SQDaoqJ/oLmo5WaTSbIkRbZs+3BXKSyj3v33w6s6mdzLoTJkQS/U9N3Z2DVCqFs09Pa
OelvG6q8OY6Z3VEjCyrNUuROJ0mknDMybhKp9k9OQf9GoMsQjMZ97Ttcyr3y29yFXLcV41R6+0uO
eQlSGDfa+dAGiHWhN9M3Gpk4bwiW/T8HH2cAZHXOiQ5HUWxBu2kdjqedMzVNgAUl6vHByWrrLDnv
XYIZycBUe2I2Mc1hHhqvrWAnJu+wP5//2jEPPvR1qbcWxh1QLJm6BsQoI01hZWODssPrxLyR37NB
n5b6JZ/zDOzM7bQy/AHbKR2UquUL/1xT6ac5Wl2waDFpyxQFNm2JFyvqmLZhKLw2jafzq80wvOIW
ghDeO6RkRtbysSLnMMQW+5CQ8hNjF4Qu/U4BoHFj2UU4RnOmUzYXYCJ85FRWVwYvQXTeERB7xkw5
FJykiJCf2MGszgJQBe5Rj4H099/rlWh4Ac/PS8i+xLofeKnTyCemoW9pAz3iOMFE5gmQleaFMSGY
UxGLV86VqZw5EalI7hvjGTBlu89roWGABwE/xJuDwI5s8ZpMzlvSzmAnQAaI6H52AgNV30tsGO6j
21BDkLi5cV6QqwqGyO9qH+VMN31ypGNGKlYgqPM+3Njq/99XsguCRHK0SirZ/ql+wY2AU+bEXqm1
RbnkgWLcToRlSBcxuHFowUcgpubenKsc526Zo3wOSvwqBFkKywz4Jw5jqAL9OnELW/Np65ACev6M
l+BBlo8l4CEdqGQg0Y2zpu4GsUgYCt8lJ3mR3RFnqq6tb5BJMMS3ltWHrI884QCvQnEaHV8MMl+Z
hRh7qAroNqgdp2armA5FSIne1PJ2wJBCW88nLvke0pYxNmQCXzlwEsVZBQeVORR03LcEUxORJQBM
2isND6ORWVwxI60ihdob/iOM7p2DsCoHgzZEre766kiQPJwQF+h7rqd16d4OG2ZU7E0jRUMlHj3l
/eeX3p8rTh6Ts0JbyznOF9DG3Y2v6FFk7F2baTLSxfDiw/R3dcSb9Qq/ieh3mKfSEYTXS/WA2Cr5
nrKY6uyV/Ynh1dIprTMMIP9nYELz5CbCVyjX/a23yCtBxaTSQkdlqh5sc6WvnBLlhC4jvTxA+k3c
1fM3ZL6gBrCk83Xf3E5AEFMlqG9xlnt3s8e2wqTCjzF+qzZgR0NyMnMy0EogsGx/uR+AO7oqpbq3
BN5GbTMNYNvCYtAZIPnh+b59OtksaUYX+JF4dhwPWtX1HnpXSgQnjxWj4E9VXUBhVURZKOkZkVVO
IywZm0Ol+44+SOBumzC7beF1a6mWzJvj4HWkKsOVlKNC4ZSD6tE3UtUFybJiuow+ZE/5sebWao2y
IX30kztF5u7zuRKVsgHFU5V44KzL+Ov5JFpNrBPQZP1adlnQ+lOmgyJT6h7plDvRonc+BKuReo0A
XsNeLEjYsEzdUxjlHptThflt7wztAV8IRsTf0nLPQlosfsjSeU3c5ZlNURO8oQSLDkxyJZRlGXe2
yMCPZaTc6/00BwWJVPQOU7hBa415UJztkV+5MLAGRBWRp/E84MdCVL6XZx6kQ2sRKaQDevYoWf0Y
JO7hjlGzT7AM1jUxZzMkb1f2UFJYOg5vM/2GXaDU+dAMljTxRWIIFjlxsMgHGa7gSC441zALmRA2
q12aqdaQ4nrJ3Yn3oNfCYWs65fKtvWaQ8NVQr7BKTuHlFIlK3aiw33yLcpeYjbngi3bReP5+knLz
B386i2EBe4K6NVK4Qs2Fi43eLKaw7sWwPlNajVVWRvwtT/x9NfU8wix5iAqy61ARGNHonWOypmlo
WfBqrB6wfsVMftuXJO73Rrc0VL39V3td01K56vqaA7+Vc/3oI4sa8q4XXXtA8QY6BouNENnGP85b
vsX2DIME3ffzF/4sdcLctnSmiRlek9N7S/L+0yZnUZUL/wRCL4d2g2b1VlqnVmZZqg6GS0lBUTxI
zoxDl7cCMxz4jX8aMzHA/dVa5poT8fBQsGxMx7m5X4uY+snrQklkX1H7BsIP0NL/qy/owEs8v5Fh
RLW2NAQ4ZCgPE1SCDsiCefN0+Uspm9YaL8iaYq9R5wDQRN8vOMmDlJEIC+LBggSunExHtMUY1i2h
0IHpm74GEN2DK56hxvtP4dkZ97uX+PyuBDEv7q8/ypL9hHGhLxvHCxJ9O1o2Ksfw0PhwICn8Vs+B
2YuGykkFKYIq0wKULRRA8GttGVUE0bzm6LhA04ICnDzMg2tZZHyd8E+Q1EcipE6wh91F0PxS4uZ2
i553AdX6nabxGSsGTpqFQ3PTeh0avNozAJv/2a4SDXNphiNBkC8OuUR8HXKVlk5GvLitZFycrDio
6+f8Lg1FT4BvH4Xcqtz+8j3dsSLpXoofyemXu+p6BiyxwwqLOZtToXPdz0bvmM5NUlroeyhsNEVS
gXQXwSzDvsA69VIe+TDYlbDc51OraT3VcuHgKUZnp0A2BAGuqm1TciW/+xPd8euIaaNoUNBqtxmP
4oSbJeIDxek+O0lziPgRRzMxP/EQ/wWO6nERgXUgFlZphOVOw6p13gk5eqbs4erTonxlK4VmR7+0
8f6bcFUrPMOO0r006qN8jxnmZcXtqpTGPCkeAgkfOVANX5rAon3dW9zlDTf62fH2enSrTmsKnuT3
I06Bhv5OlHl9gqtJJl2Ws7wq0Nu5+WSK3Uat8jC2dVuyJcw3WYr1lpbFgnDn+RJ4cu/pIjr5qf0f
r6v3UV+Jm96bTh7Rrav7mBA2kABSEKVjT0lRr30C9vMWLtRvEbg2PNGlU5bbiBAmh1qkIGAk2MZd
VnWDvL8WElnBBVgtNKZs5uLwnO7A0ZUyxjVLA9vDAljY0K21MhEk6YesJLlkE/7q9bUlhGY8vvlm
2erDkyTHNirLa4xEL+0sy6lI3cXjOr41c3B3ZyVmH1qiOeVssEZH4a32g2rmB8LW7+V+zxJbjT71
HBqo/mo00Zwi10rFFOZivt1slrBlb2ylV9roSmc7Ws04qQTRjLia4HveZratunPCEqMpryJrZgZM
JyGGtC059Z89rZCMd3Pq3NT+JWKapR8RQwFi+phwafvshuaFVxOLzoe1DakN884lzP0lxAOPD5LZ
cFy10/PDYKhPSSmrNjL7uXnWu+VtBUhT+ryG5dfy7ovvRZ6T/32QOjqLvhPIUGEY3RlJS0eJNHkp
9GLjI2/2xIwifbHaxJ4fPG3EIOjscGpcKtxAjSIAGiFUVNfwj6SBQwak60xRtpf85PjGLgAQd7yF
mMG5xO6bBVo9tUAyLlHoVaA4ZfNtdbXobGbfQjT+DgvR/rWaL92q3/S//N8BhhuojtrDQnqHgqfX
Q5NuUUJlfYg9AhaaIEecZM0d8J1ELVAlB6zSvTGYviexdN1Dudv09il+UqWopk/Q+wJHrR/m9mdn
Q5txcbKaEpwBTyqzlq7CyiMDzOHiah86mXG8OL8nmnYRDscWR7ujJDWLg6gFKPmEHDIw+n6UHjxa
pG1VD93bgDHNZVa8qcuYzSFRx1M0T6MjeL6puDbIE5OZf/MeqfsPqx+c0y6W3hr3rLp7ZeHmgVMz
ANTc4E7OTGNlZs/n57qHzss0x3qOwCAxeV37fiL6aZ4QP7/bJu5mPII4GHB5LY95VKWwAGLnkYCf
5z2Lu3gfvDTAfT72b7TydIGQuGjZqWk5DIPtzBoWhUYhNoYQVJMk0bJ9UKbNUyUeKEVQuuFywjm+
aOeV9ly+KtqzY0kX/M5vUva3ERQurHvODq1ZuLdPm0sEQhe4oJBYP47FGm1w7yoDgFWJkLjaSnQJ
HD9JhjKgpeOduuZgmwwZ8aFKyX3vnm/CvgLt1EjsKELQIOtyD5fHobtTVY72DxmZzA8YTiyd3dOM
GV9ucXgCwscAEyMzlTVO4f/prJGZj5wJpbQxjV9xpUkB+ikSHkMgGb6Q59koY3D7SmvvEF0ysBsl
/cSMoq8TN210uaphlVZU8gJRh7NOCCdl/1h+YQ0muy74iXoTKXGfPwIDk2FXPg+EFKDlN0kq01U8
g2r4gDgylQXQqPITehBlqu+dg6erM/yQmfpFIqNB9mhJCuTUsb1vj6BMrFrT/5gizSnnQWQbhQsA
3My2ft0EwOenk/ltA6atWapmwpRAWKE6unV0nCyg4OCgoiqyQw7WK3/I3i0hyvZHD6MpaZVw0ePt
7vpVL1VxAo+GYpMp5JTi87kdBRM6I0mFuXKlCJJ4NH2RZ1eERSSa8R84R7el/5eMbdZ+6iTvY2nl
UvxIyWt9Ay5bkgoJR1YcKiDIuBSEMGEZvZH1rz9RmDbNe1qCpDRsxAz3yYVQg3gYvMXfmsZeEr+J
LNxF7nL/FqAWugDwqiRqSVPO+SArlk3huyCCuOoH7EAkuF1JRM5ycRel+53xshu4sK5oxoiTmk/N
SrqsWuKOjB4QwdpI213HpKbExiqUZg+K5gCBOIaQZXpdOYYKgDgGMjvt7ioTHblcxeUvXpxcjzqs
T5YbvnEf1OCHijLYStEGDt3jkLqOPrDpti7GUmAwoPD4p2yHuF4Kvi+8YKEKLqMkvTr9xpiuCVKz
1LXpbT071tBsqxRXPbc8KHACwwRZuOXK02GeJ3UPue53TmkkKPBsJ1K3IIjaMl/oCQ/PSTb8nQrt
1ZbQYsE35YJrdSGoHgi/toGmZfDJRiXb9CODxWdFIPXY3ApksCo1wlwwVZcHQIqcmHb1xoKxy/S8
MY8Dy0OD3m2gSRApxkKzg/9Ca7sYv5TNFb4XQxerOrElD1G3hasXqUTNOVkScJQ8nJueTglszz+m
MZjMoui+am/fcV+qtNiZcURyZHpGurlPquU+ou41PCpPGVvwUH+hGpNOYjf6uzU6lQRunghjG4ko
3DBh8UubZsbQYRJS+SDUN64mNsVbu0ZV4vecNS6nZxnY5rE1uq3pLjU9lo65McakbYewWp7UXV6/
I1jtv4Zyafhupd0yWEzvMMR2OCAF+fIS+sHHb8i2mIFEaHeAp7/5bj8/gIVK7m27gDf60wHgz7Am
TSnpZSIkb/b9Ydc5E7nXOUfsSvkdGO1IQmJDw4dUmwCQ5Xy5C0d0J2Ozeh8Aq1h0VAW+jmCxHa5H
OIbB+WVi6gT4vBpL3XoIt+U00/q4aXn+deTzixqPZd4o0YG5Sp6JHKOp9TLI9f8VZm+nsWBeoZpV
5IuEjsRsKi6+VeHdxxtYhj6nJ1eSBus23rb84+UvxsWsSJYSNus2VxJW5IgSJBZiZjGxu5/tWv5e
a+OJJU+TexomePe2L2BpDvpnMLnGFUy11qjRjP2bldLWr47GsCLmgwinobpOHaUraSqx4XwWzRkl
YnHENpIGV+AG9Guh0lpF8vvK6PMNfQ16xXsjAr/Sy5RYozHD63WeytTEhLP8YbhFbrADBR9jkZoQ
KP+8QBrWEYV7Kiq5DMPo8S6EKdWRZWvKswoyxz0jpNhtCjQXapWdI6MVEf2rA8N5UmpSggaWnp0/
+jHiePK8TsMKXVoy+nhOgHSRTlGrrsA4IGuPniIepRvA2KzfmhxnGosuB77nPtWxsHjzTAydRWrY
q15t5jkoDq94nCJ+v0ZfNTVsg0Mdxp6e94QO9aEw8hpM/welR07B2T3coEDV51UnlZlLqt8oepgo
tG2EFHuCSgumc9ttW9E/6DYX2wOdcDuEj6vpHwVgL4TGEwJHq7GVPja2f7A2tdekGxzzMSrdpDd2
YYB3Yg6yP2ZtIcEVBsBZRMDuTFH9FPBsh+93R31tFcefM2XjrXkZkIiLfWUJuzpcOCoCoZDopK9P
i5YteGMJSrXRgVZVTPoTCZfl1Mf7VU5jSXwqUYI6Q/vPiyHJC3KI+RgagbxTFwf+dwLFHsgVffVM
z6BkADZ2T8nFhsfjIPuTxDf668r3QhdodqpBSR3Vi+tm518mUOCZxpkW//U9+ShzhVxREe4pn3YK
M45OS15Dul03eQSP6trP/yKtVFYp3D+BMyl0EGgQtncZVzy0Ins5vYxrW84pAso8z6V966qHuiGZ
b1tb5p0QaKJruBjOaR7YOdquso94HKEfrPmgOr78MZTvoxicfLoE7dFt1hzh3QbeKG0gqjLaKkKa
6tiPITz6iw2wr83s6KqpgILymgLnkJHm7TeE5tDOltF1S9qEyC0dCzC76HxdhLt/5qWqwK48h7Bq
WGErbITy3hZxg0LZWj5AmGUYCYpqcjnw92pHyVDM+LDp+XFP/Yh2G59NsSTa1DR9HjWi93ZyWc8P
BvIAHz3ZS15fr2fga7mFWApfP1Uf/TPvPV/W+vcBrWVPPqGvUnxbueD38j21XbywDk6joAmWntXF
0Fc9KE+WipQwRJL+iiv4MzEnY0BX6DrawCYJCEAQVaWLK9KfUj6I/RVTRwrV81VFFkkzeJLdrZVM
yYAOBrToxvrGX9uZiXzyQGAJk4vKQ0UdhvKVRzaT4XyHSggqGYBRpRMocj0lSFEnXTO09LzmEmbx
HbYvMEFaQ3IL2TS4eTxk1g0nsys+AiO5g/09/ffBcdaf1AiYzAsAV1boA7wZEB2lH0tkzMwBmeuT
9HG9SlO7N2hseP2ye+ds864l5ppQQIV/q5y+HG1nttrgKS5n76W4T6pPoE53umcDyMiqyDUVQNOu
qXABpzSjmihy9uSRjnHa6yWhiWVh0eDhC3QByirY7ERkpCwszvbwlTIBhmET3qjlZwLwHn7+1K+9
9bN52z4Y1AQrvzegJanRT1M+D/OajYj6lUBbuZawFpoudhMuA2H3BalRzxeU45XgyUC8AhhGymRI
571JY9p/SRmNw/AXnx9CJWUR15uo05OgxjNusTcpzxQRzNamwx82aiIY+nyOSBFi1T2wzHtoAe1f
5EfGb1DuLD7a3nqMF6+0hfnvC9rwVq0CeNuSqvHBL8s2tA67MKqd8+3eA0fqaQfnQExJokQOKOu3
Jbgh0eYop1ixME/XBbF0kyKyeIR73Ixsdjckj6GhuhuEOhuG0D3l6ToJE/08Osl1AnKlmRkHmXS5
+8BIXvzi4La3AfsrM9if8P4TtPG10z8j+yhUxUlzJwn+88yagc/+EcvAHXMbejr/IKr5nurMpuSE
R63NAry7DecEpT26LvQ0Z6xn0SR83ZTBTfL1ydOH1aXC6yJ7R0MjhdTCfyDHQc9ao3QGaS3uZw+L
208sxVBCRjYyMdvJghiOIABa368VveFDmwJi8oBxMiXHZEtffLZYlq32NdwSHioXg96xrXB8Gfs0
tAaN0463k7QpDNEiQ/iupFGJ5/fl1eRBztsYJdAuXIe1oDtUOPxjSeCii3Ys9Gl1nWaQKo44Qbd7
RLkC3aoCBsPqNXZZdePvvqBLLD3cl6khGw4eBPpJg4UGmeigJvX/EWP3RF9ofNgBBUiXKDqy93s/
5ygb5fm8ujV5GsXgfCVUKgMcVIqH4y0nmw8lWiOpFq0wX7onw9FNxKzFndY8MBNaOGOOPnDUi2Y8
Np/400jUpuS4LjqACmdVnS0u293uQKLCCTyb9wD5+s5SOoG+YjlpJK52wfhkUiFvU1kmzoiSC0PA
mvZnrIaJXoIDiPhOmp7FiP+i+V7RQ53cI3URyhg4lrR0vyVWsscn7NztCOSnL9V4dz1gf0CWs0TW
6DdBSfpLoTIF1OxOwth/fTgjpF/ZyB5UeQGirL51oJqZ7LXAaOkVbRzN7r2qXRrKGQLtOj1rOsyX
9XTouK4gkFpbof5ME5yvd1uCHgDtjQTFOmOFhUd26/iP3q8maVbCduwpMjGifQF4JLmy8HsOYhLo
D96kn2Ih3ZMBgVyK0Z46aJjm+659JCkOx2NmAnS0Exvr4V63cu68rky7V9iW91Yqno7kZKSBR/Pt
zuOeLSNXpuhktmfnNuD50Og+tz3Wic7ywuERJrREkzLthfe4eSoT+tuO7gIAftZ5sO1Vu20HnEr8
nu9WeTL0pmLODZSYc40fmbh2/YCe4GZi3zGgCV/d09xpzwikB7CZmzFHWYH2tYjsSbqyDk0ARgZX
NbwYI+120Q5yQ+tgc+UNNMmUJ1R4gCk7or4wb4m+8iq/bjEeb/vY86z7iG4E61u4mymjR7Y9xh0/
AyFkLqcrI8XQCtmdKCxfVJdd/mpmzMhjheDro1e/d+56Nj6TMtQOoISPVpfZN5Wa/1SjvumlCWxw
3SxkEzQgljl1bjHVGs7a/LqK7CgDaX90gLfBpU/CrsXde9ga+ld5DKbhgTRC8zTYpOTq+7yAnexu
ZDWyRG5MLErfRY885+5Qj0QdO+BNOlBNDgbuAf5C8XePFbAZ9FbTFoHC01hZ9X6CebD3A8inHSXx
Gp0RwMRdJSGywsyKh77rTtRLg3CvYwN6D1qJdxEtQPjiniNtcVUOKjcAPlN44Me8ZqqGv9stpa8N
aaoE4JcNu3jzn9vznr30fy2eFAIogGFnf4jUbQi+2CWFjiUJeWcV2gRKwQDJwGh/tDQDSjsmOQ6V
HgWYDUU1w11DGxMn4FJAniXfqhNni2Giy4wKwyD0q3e6Nv+0HWKRrerAwfF4XA6d5BCsSE6W3XwF
WpqGRsDRIfCg2FjKhil44+ZdQh9iJ+lYQyozotQSfNxp0lMosjJf+t59Yv7bG3W7OXpdXbF641D8
mRgDbTINUnDpxfunO6dgIBI0arT9S96I9EwD9Q3yxNpScjE3/jLNdeLWsislM/6QOhNK8NtJBbYk
pa1TUqN2iLCrusGnlIeA90LBzxJa/NHGjvR6pyRkjqs3qPlqePlfWnSOmDXAft1kUX0xASxRg2VP
Ia7zBMHFmPOgZsALb2tQg3OMqVcq4dxIuHUWOvm9vK5TApPBzZHIu24v1LoCQZPqWsYVLgIT02ER
xa0BiTl11p9zGOMdnTgL7z0dKZE2lOUDF6QI4+9vooq+ekJoWhib8/GzY6heakHsaPL4tpVFwdzr
zTeKAWMqoEjEgIYxPt0zkpOYHsbx5EqgobTNjrWK3mscFEARn6BwJRf0vEY6VbbIPhYedblt73r2
dNzdCKYBjAIdEujtKCvHGdBjPyJezSf3TxinDPtRB6AdfvRe7uInXD4RgQhTW81edoG/K8hCIDwG
7UNL+SQb4nhS50s9cQNU9eFMHUYl8yo1bWNYECWjUQEw6kKZZdtpy+C0VfeJ2eUHd1u4lZwzsraz
SOwrXKWLKBreCbZ3c1tPnYRpfHdYlzVhUh3o5/dAtwM9jOz1Gvzd1ZksV7iAxmqlkuqO0tMAQbqg
z7ZHyndxMzDblvoXbnO9ndXmETMFDmMiHykRw9MVko92xbXB4qzb42yS5N4d4X5gYgaG7+qeyjUv
xMVAJsmdVwdJOe/I99FB8E/2K17vfZFof9FBQCvhBqXlJNaVbzCYJin73SRsSEuNBnNr4Ja0ACcs
aduI78lxivGPqmejp+HFG2fxrqUFFkMYi6trc3w56sY/cIdfPqysT/PowSY0+MvVQfC4PHC7aJRb
50pHrpPdftBvje5MyENVPhIFZF3IR4tA+Im8W6IYNnlJpi0iTC7z57OWplw5E6RjfA8NMBO683OZ
GRkLgXSDt0k3yHNWSPPaDSpRsxYD99ansSVLgaJeDAVpKu3PqS4R2wp9sIEkreIrUHcXEEIMuCkN
qMK93EBM0IxYJpzjc/yngrUHK+788pJryD2WNYl5FQ8tP2FCfDUksaAvo3OkcvyVgoXROBTQVI5O
2yGXIjAO1Mks3wL7vPSpkJ1aTHDALSC2//lt7lpDkOiFKJU/NpeGGFeTc02BOXsKh8tZnHqQwe2j
fEKkJ6zK7k++VmT2qbbbdsGxTnyspQW9RirAP6ja6PiSB1ysY+GNFqltSc6KQtKTAlKS9VejrbNy
UoioDzkgAVN9tMrpBXh+qrTHBa7sUmFSIhem7Tate/j6fluwBkMi7mWNXMgu8NUh9rgtJsuISUx7
2cXTqwbp4un/tIt+1/gZ/jMBM03GWKlOx7ILjyNOitl7EmXlfD3HsZrdqabX2386Ac283WJFsyI9
XkgQqEM/Jr5nUOU3F6ZaSugJB3gp0RsVeQuM4qNjj1zqeNM6+ybMEbE3aQnlwLpPA5J5iwMzmu/b
Vompo9mKvN0iu3PZCoesIvw2GEgQWRiiCsCPhLRax5RyYPdOYmm3h14X9zYov4a2/nTXQCc4ar51
oHEu5V9Of5mnVi/oG4SBkpWk+nCHn/UxmD/t8W/f4JtitqAIZA+I0f8wYZ6D0BJ9KIb3LHo1AAyu
9L3IEy15B4FtGe9uR8P3s2vd3VkaKZjFwXtz174OWeY0s8DP51CYbZqb6kKdlUIHR514Ttv+FcAY
Lk1AdiLwDE/S5f30FA+rCvVLgQir/DbkCi19PMPxm9GcHWc2hck5MAEaBsdktoGNdOY/H5DxcdZv
AwLOJndiriaCG7koT2wAd3GX+A2rP0xw7tYxQjlkvcM3g8fMLx7xTUkzEGQa3ixQnWcJrZSbkHFU
6mvqB2uzOKWyjHGt5AZ9/iuVMksf7mbvoD8wWeAOx9t3E1Ma52yWj2eyCMCoxUS6LPCzfEK5RufR
szWr1l9g3fow4tUTHlC0FxTtjE5N94bnFaCvdjb4bvfExPbBB0KG5nGCME+pMXfOxptgcCJsgFaW
fVz3LN7EHceUbVuUIlqTWEeZg1osNC4iqDjOG10nrcyBpnMIlqOoU3eXuXrSEenJRuqOJs4n+/lT
oa1gNC2JV45O54hgfogDM5pZ65awy4EWNaCgjzjfanKV2uLW+4rnxwGNWzJab6saJs9dlGhflwKE
A1bdzXe10sWf1rVPJJEuxWxT5fqvRxUl4CH5B52nWZfI6kIIg0rX3k2M6+6xTc0JAJeZSYV19zt0
u0u0ys8W0SkbDVe7JFS6P0xkhyiHEtBkcBuXBpyXDUt4X9jublhY2oWRXifU8qHueBbOfEJKUlo5
aeR5uJ53R9nuCrPo1s71oJOayh3/YH3dn+Kgz2Jq7Ud4XfkcAiOS7mETA4ZI7LWe9RM5XjSDog58
BPZQQNtV26u36T83j1bxKeMlKMqbSNoI7CZ1r9UNHEjmXDBpJLJI0YGsWWKtnlkPOj806PeEfyms
V2fldC+38wNU4gKg+ZnFis6nWCbEQjbBS1CJJn2CClDsEVim17+CmSnlnKsGQIvbzUVOtHC6aKAI
tifvEkUJRR0IwM3xsZLNHTmaFEz/FxQKtTMsfikmkMaeJ+duiDcy9RPiU2xj4rHNoKV3Fy+NXgar
1esAqu6JyKqFtI7PIyHCiT3KPsjc6GdFORO9uECXhIOeKTV2SuIoy9WVww/KXvxE+gI/JYyTLlqQ
S5G2Ogqf+zVISkfYp+KEXlu3NUnLaKqnnwJbo50RrIiNGEP3ppCsT8lnFzQJrQeg08iyzoZ8ptqf
DPT1quE/Ar960ED7PNScL7QjCeTo8C7Vq0biyPpT1SbC8mh6uSZKOTspaNVq6k+zjclDIfWwJBM6
n6Zrhl4x2qiUsrh2bR9VvdKKbLjaFVJ2A4eG4cNAP2zDxgDTgCaejskQWE+NZ1wPDuaY/vQ8HEXz
zTiZyacLViR4BYrXgzJkvzSGkE+0Nl2kU8We1pCbPs1fbET51eIJBnsvR3XnbdJBcbOU6Q/FwUNJ
2hrPpJmY6ZAC7TS68VLkZZy3Wv310atrFz7iPaMBd0dA6Zc7q875tygoztSS1i3Rf+uGI5N/0EOq
2gWrifyCx0jOBXVwkZEO3xE7yKauNf1Mi7LE/M7zfZGkyxEvPJ/HKcEctMgUmfGBoWvNNNjzl9ur
cxTR5hp3nOv+L1SZM0uh0V7QjOeE+l3478PwRC367bsLKMi1SvopTIDM4rmtLnzk44cyQKRFEz0i
sWhkUPJ85fh4ZBLqGehW424Fq4Ibt99Ej2CNTYJunYH4lwUBz97+t3x53G48GAvC8iU3ws5Lstaw
pReSdBsIed7yQtgmeRv4BHcog8I79XqXsFOeVijQIX+8mC7FR87u5Kis+oB6D40oV6yePoxZ0doK
5y4bi4hIOCdPej1q444ZPDbV3b7Nnfy4Cvsc86HBOOxSKD9NjIgd6bisLne/yN9pp25Xxv2up0Z1
Za7jfEhwgawWCMcR2dcS0auoNM0z+JgNB/dbgRpoKdXnXh+0QaOzGI2tseThBlaYPo4mIMXM8X7e
HNb2ppUNK/pE8Rc5K+9l6Xs0Cqm8O0aFht+MWWLXt+5jtkHTOLkCOlfh3iuoYJ8HyM5MBKnjTdMs
99ywFb5bLjs5o6ELL6hvUufkMKL5bICIqh8Z2XcNqUTUpq9ChNjZfJhiUcTyoWYYZW/bAGsAWuWK
3GTDP+jEJBx+U3mjYS90YlkBlOI3Uvcvxn3eT+PgdTclCREHroQDdTYrwDLcW1eEhLacjZHjNcGo
/ySh6rTNUNLQSh5LjQkjmOp/osEvq8+cFnqnMlWfVkJtT3lKiyJKeugxoZ1jQ3f2aWlx+q+h04/5
ftl6PkfgLHj6+/+CDZ1TVEt/gR6JPrFthvfiG9yzWTe0jJPFBRoPASpLLtwu2znKwxpcPCFSyVQz
UxPs/yBAEhfzSYNt/OmAorqEArpXYM1/VLTqeZNpt11SyiHGtKY7er5K9xkRuySoGzJhsaPHeKcK
TNMRZRtMuFtJssPIANJaKmnLF6pwdx4O89cauW5/cuFk3CLZ6oCDr9NbGy2NXvdwufMGmtwHtiIE
GhBwMLX01hCk8nSY3quvPCdjG2BlR/XqTylYssdK4fPEZRiwaUGy73i9RvSqmmiShSfp3GGQWqh6
CNi6x4bhvGnoAbb4vNGMQeE4LOQJNdQ+1GJ4/YHR/h60ksJrKR2s82ByQuYAEDNpQy2qhG/fbJVv
re32ueRVyat3dTRCyMnnjBTp3gsKSHjGycFa5/WCE2e4eGgb6LZiVUXDZdnOWG81E+5ZzCGc3Pv/
zbDpxjm8uKlSyhWLrXZUQ/XRHZGt8NnM2/q+3IyObd3m5hguLWe04gPvV9ekTxM4vm78aRkP2IAA
Z8Q0MdZIgUXRHAsp7HzelEP2Lw0/16cZptrRXk8Pt1BShe7ksPTR5BdYFx97U0Q4CWN1TRo+MEpP
GuMWbwuA8I5tGPBwat+ObVze8+LKPSOHE3MULP9/rN2ZmXvwz0hGHxKWC34tzz99kkGWZzQLrxRL
OUImXE2IfaDjWiZ8HFVSLKkwod5bNrebY9EHryVYpsZ92andGT2X0SytX2B3mW11DCLe/XGCzyxQ
6mPwm0Du2c/rbTSdlxeEMNhHNhC+JnwyKBy/9miVNDJ3SeIxU0RLcSrHa6o3grNYgjKgpzn5FhP0
LG/4sRzBsccuc0nbh6VuDn31ScM7VyNuraTzPxNPslBgOOGfFqA0JgBc/S5W988Ha2dCR1o73lZr
0VV53KiOHroPT/n7Tj9LQO88H+luahA43UF1Cvy3XB6SFmJaFQeQbAaO31Qpu9hB+AndzaQJnEc0
oQ3WT5quHGzWxYfj9W+x5oUA/cUoPRgD3D59YugJ+tLpdP1giqtfTpmpIVjVU7gOiIXDqnPNOFtH
5eCNwjHAjm44JnHL+6sXi3+l53cuQvjkCsMFQOPnXsebb48Ye1KuHukph/1csRRDryvW2iJgIDRv
hEx7QvPu/gwpO9MTL8CB0RvwWE9dvT/VTCshJlafB8RfvBUbkWtdsxGJlxIvEt5/JI1d9NWvf33r
G1/eXqD22dvUnA4WSeIM5inJre2zgGPcG0GcJe8R96WsapoVsdLMfxy7C4zawW3UVSqOVYndKM1J
QQsABOjZVlVdMZJkekta8rEOKRZh1SJVC6N40vZq9VFcOAh3aG+R2AXFHg2o7JRKekb+gP4k63sx
3/zfmIpOjprmlLXXXkua3ZBfPcQ0aPQxFkpFmPI5M+h4tdL0N9oXTqB2QOxOKP7Gaz3XjOwKo02G
RGk/H3gRgyA/RiB0q6JhcMuAstniUixt25eQm0f+mtF7NfNlQjn+frkVFpph3Oi1DRBxGp5UeBmm
V6Xo6/gVfTcFvzb9WvZY1gdHuIv5qdAh2REVceDweH1WMzMx2Pse6McB/feQtHR01QZhFTdrOpSJ
hh29ikwRHgS+UbOX7AgmQTEO07addNkw5uuLxL/F8fg4Ipc9E56yX9YGf2Ym7GgDw2/D0aLCWxhk
HC+0evpmd8FqlM7XPxIAw+6U1l/z9uft/sUZqhigZsjFjh+K/vPdGiV8Pu4IRIVK0gK4/OOe+GhQ
2iVAxuddLZBeRQW0KB39D9Q1KdScNNdA7kuoUQZSD1PI7p/8pu5XhlWZ8T5kzai2fV8yhAuI2lvk
FSXB/aHQLOvQepC5QlDyM1trfh6V9QRK1MmmPCLgXU0a183aur/DOWnHBVItnOpmlHgZoq9jgCx/
8/56+mwlEzHKkXdbsJVDqWd3oGK6Uz4rIel44MF2pAH8bU+gw+BGD8OPMcLDylPTFyOYSzIQylos
7Njh98ZVs0mPmF7ZtO4AvbkUHBcgujhNeWNmyt+3Z5LJXiTAAPA11xH2G6111kS52rtTnx0qKcd/
KPlULlWAKwmfc01DVCr3osx/PuokeEx2LGB5u8Wr857tK4GWY9JLA4UsTr/Ph20K0oPs3Koy9yUL
bEMDD4L3TM0Ewex1yl6/i/R3C+7l6btEWDMsJK3ptdgV1p0Ls4yy2wAlS4bHGKz7bMTf5/jpoM6v
Myyf2KNfesGU8Gr2eU0CK3YrNOS1eLyjYuC12lGaabL0tpU8pJ5ZN8Yu21BIaPLW/BqLIOPiH3Sp
qJNIqECg8DY9zafW+32uIlU89M9hBDakqzonA3/jagRqlWxUZTu1d1nDXqLmcyQfzB5K/jwnEWWP
LIChRtU7xX3IW57eBweD4pHEhGIyV+Zy9UZykRbildtB9/vOuYgY2WOZqWkJSmV/E/aFcO+F78CT
P+HNTu/MDdYhM0kggapMKKGI9TkHZSeRg/6p9a1ea5eGeKmNfjpydvL1wk7qP/Hi+7XCjeyhBthl
ktCQ+3nbf3d1Cu3OTtLoDISG9oxhUN7D3NaW522j84PydbSAy7PAjyYorjcXkqMnOnrYrn8BJod7
VzZQVUz7NqYsM+sx0WVYBCXT7cpj78E2phWuuA370l5zW17xHhyZMTXw3jmDk3zLGQuowovYvcvI
7uwTAQl7AHQq+wYbR/JzXa4wkRwH0vEKvSzAxM1lDvHY7E1KzbIvBkZCtCRUIq0s1BP4ufL1Ae2i
V4pap41CsKcpXZMLjRNIYpIZh3OWXT2Fj9dbYc2OJgCnfZ8Wm2aJI/HkHOLVUK0vv8x32/Xlp46y
KMOkGrfkb3w9+Ifdlk46KXRbQDJxXIszPp/f4PsD2kkBbF6GLtyIyTs07mLWZ+XVWuIgyzT1Q/hb
5kPkOB2g9Mjl06LIkraGq9iF+1cFF1KI8RjDL8JymwNhqs75fbte+aoL4lJx2uAEFyLUrvkuLu9g
JHpqGnoxVMJxQe3Us4EQjv+6DtOdpAYNz3v25YAU7ot9sDKhUGOXwSY7TQ2zpubXc/QzahsetZJg
m6DW7TkRXS/kvP1YEMo/vdA+g8sSmcI5bh32PLiN5LRTA42DKMyYhGerbPUeCLVcSlvivtds8YOy
6dw6PvdatVrXpUdkieznbBF5gsEtu64NXAYBKWVoB6RPAjjYoXgorIGnpLf3PulUUKk5Wb3C4SX7
glEwYO/pkhmYgn6SbDbnKjbdflFU2Y+5keTtxcfOVNBHWPh6iUt6W7Ow4ZchV6agBvahRF6+RZja
HAuxG058cVre7TMv6xrOqzQp0XO2ggcdWasw3vB4cElcwi0BLAKFlc8BQN1qulxvJJy6+oHmSrXs
h/Mqd2p8/Nlb3wWM43U8jD3ZB3Wl8bWs0x93+bH28OkDIRjL6QtJU4iZ/ch0FRDS1d9auaBMej03
VRMHVFsbiC1Y2SEQwrwU6iP0TG+S5PcEYzUNi4jMTHsKdoxZOr3Z5uW/ecwwTYQTYiM8ZpLs7Vz2
QhdAjNTF3sCcDw4SQDWHgp0fskp/o64t7NuAoko+DiEeM6M6up2m0IIhirlfeGtOB3qYd5BxfZiT
8MBKYUHNUjKY5ULrQNga5eO3trKXibVBQyNvaEHruPQYiZlbDa/aqVKmtj3agD7zPt1FOrfREEov
y6a26cD43/McGMHzFGHCSBHbuQQkJhIQU0gmk/ujvlwjDTvrCgPTr4cmh7yPhxJ+ILrrleWcq0Em
mfvtnqxhj2jIG9qqDNwbOZjyDVL03Pb4Xo7Ky5y8aPTOnPofZ9mXH1cVmQEfOysxvnx//xxlqT4q
BIGcebiDSEgU4q08AD7kEYw5A2Dwr9cWTnzTDNR6WvMOOeKPg+J4nXV/kIAvZZWCzHha5ySePm9s
+c4nja88B4JWhaU3y09ZuZI2DRNlD4WIREYMjoaYL/BFV6zUVrJlFtc1dtfAy+Nls46ITSYI2OPm
dMtZdZVzbQhUokNxG1GRwoj3rdRxkGk8q9IBWHnA/sgEyVw9mrO6Y7BlK17hbNKdi4N5KOw50eyA
bnJtWm20EldZ/gHbCk0eaSkamA7gyaogFzfM81O2tcoGl1hZuJye3FPG5YLERtHz3NTp1des+69Q
HZCuvTUwu8aWr0c/vGXol7eJAOKWqNv98xMyxDfFygGGHUYRw04azO1TJeZZjP50aPwKcHmi6aLY
PKhm1COaZvLG+13KIhxRMWHA+eC1/Pcqh4P0aPTPYo7PilkLqGVI1dirzTV4JRQ/P7JIrdbOST8X
Vc/IPituogBcxpqmClSMXSGZT9d8AGKm08OU5rWdWi0YdOvVlgvEMO5ezGjisRleawx1n/9uAtaj
Aced1A02rhv/dbDlhhebOBHRQkc2L9zBkdprL2oSrY28piTEeKHaiVNtZWgD6yuBDha7gOYgmRS9
mWHY/NMYln5F6icRW4HRgdhlTMKdYaPkTNUCDe7h4qikaUUkXRh/jl8fcFfnu1RXjOFY7YN9QZ5o
CGRov2OuQQZAwEtyT0framwDH5Hl/LKO/bceMGsxP34lllQ/TpCuN2moO+obkMZcn8zho+LWzrJ6
xbGbF50vg/AOusD1PGrT+0HQwy95yYNXj0MF66o+/M/zDemgvIJYEAW3T5CwIw+sCzONxpJ/fxfU
LcEN/WFoPJpmx647tnQ9mp/Lf2UYLOlMOzqQdil4MpAprwuq119jL8BwwaZEw+cxeKUGYEDV5Drm
KmjKXbkIbrXLotEv8YKRZ3v+kpRFLIk1IpNUkZxAMad/oy7czYwEKGFOPplMFmq6I+/Trd+QxFDa
MrbbhI1l+CWjfvWKJwEqwLjWGvyt0ekVsAomajMSDXkeGzT6A6zNFtA6+yyXozw0NElUvMmwi/O5
dEVj2Fp05K3qKz93juHzz3YWp6VFPrq4YJ/ShgfjMqTqlIszUMy7R1S6C9iDNX3Fvvnqdm4Y7rKW
BRL7Ya/x+2WufNbttZyO7le+Tt8atpPelh8aCOdAu4Xyq9npbNFCIBdw0iZcMnZf9S/qZPEIZeHK
UNXqU/leMplkiUC+DwZNmZYPqcNTHT6VWjl8/mILKJMD0qfXd2Q1FMf1HQDp9QIiD1/lyHTFNBSp
oFyl41aWNxVH9ErBtjvZXUm2m+cGEdfjshoERLxikp74FsP/R8zFcN3SiVUE/3AY2h7+IUnAQrRk
VkpiLMw/pViMRFSUZcPUqNmcQ0y/8UQHxnTMmgghO4MoEajHkV9R3oAUaiIZ+OGxiz4ucoZDtztx
BZMHQEE950PPn/c7x29v90ndQTQeZMx5vbSEZ6FvhH65eQqDPX7/2DpEmtl5Tu0kHA1T3f4FW9/w
8xGn10O3VLAwCPreOQfqAoHGFbdAvIGV02R6IMJDd9KyIhYvjaSLm/w5hGDOnj0CV5Qk1OAZI51i
OYhiYeiNteGT+7kO27RxjSMROwtCP3CEaY02+NxIUtnKi1zhx9Qs1tzpOT8vXJOUgx8zWKjmoKXN
PqaKNR0Be2B91BPvRmz0eyhD5r24rq7PRtMQaH+BcrtB7evRh1N2/X0MIFRNlIwgMOF+kLhhpJMv
kVpqIOT9xJMnsPTLiRqbEIpt3qct5S8tlnFszeyYcp/dC5xNfdl4v+7WzWQvKahHt1p+Df5Ag80M
CPM+dGLjBW+qkv5YrGofBWAeun3dkbTzLyV/QZoBvEoi7H1eFuax8KC0q1F37xZN2N/C9kUBTNyQ
XCPrNT9uRlGYZLXgfiiWMjR40pDxhzER15Sk0ckGNMtE67v8aUjqXl75Ed9QWOhEHFPPuZip/07V
0nBgd/Tmhyo+sOBJUGNwsZ4/ahuxak/jS0/z0Nm3GZbRJVSoIqj0cgQDIepT7T9jVDX9S7ReRaBc
CD8ynzQnV7+prYgRCRPcLJbnWA6AP7I6pBtYYP4Q4n/W1fUEuGgXrQ1yvPDZCRdo/bBI6T/HbT5s
sRg6MpWN4kTindhQ+/YwaycPbLVmY4W3eIvLly+NOwcjl+r8uKeKoXt8B7TcYQp1tFWYexrxox2f
TGeHf43iK2GiHIC3/pyoAxnbkQ2ktndT4q8HUKsQBLQo/u00XuYkr3j5Ft6n/cC2OUiFzgXBfHmP
Ee6c9tC+hRO3PzPslHk9YisKAOzWeLDSUB93qsyMppGCM6w1cOkS9c715utjlKlZKB531Aq/fK9T
TknESQs9thMRBvRTXW8DVg3vQSVi4G5BB09tMXLgG+bNRbcanqn20Xq6E+PUwj0S/w1DG14bwry/
/Jfw4/AXkSaFTACzAFgog5MqhcCB5kYfDH/JHx8l8SAE8262xKMuPfT4HgPA8tXuOgNwmTgcyMTL
9P8Qs+9YcaHxZ+8lGAo3+mfb00O6lYfT4hRf3JsuG9lsKLhm6A8SoW/7b7ycLxPwxAfFiprFH89d
+u+LHL8dvgtZtVv0iEceb/I0cBNmmqzS+y3i7k0002dW7gXQyc8HFKE81+v923Ia8ueltKVvy9uO
LgKFxKql2nPgeC+AVsxFiLo9JryL8PW+YnnU8HMzj70wlSIWV3QdX7TIP6mhMdOxDeZlSzsYpXf5
Pjspo4gFJNpzARkjci4XNtlBosRcC2zuVrB3pZ4zdafUbBxiDI6ZHTYUx78KcvrOZcpvIp5j7QdD
51YohLwgVdTL+BKwqrkNXCthg1/FuIl93kCxqtoYs3yTgB7AGl7LBfJPY7nGbomuNN+jQF6wKMVJ
jPiDEJeCM/TXJhouPyXonsS38xyzJlkZgt672HV9QX1lxVOf8H4dGm2jHXUddXL+uJHdlVtyj1Pr
Q4uaMEU/g6/SY+pN7xdy37sv13W/kRU51TWI1UZsujHJuAwyZdzsChjVwh9VDVq32t6LNghEDEWN
RWrH8sHg+Yfz3XYHdhwBzCp64mJfSWxVOu4Cz/TYZXQ5WtGDQJiL2XXVGU9x8uzF8mlgz6C4I1y6
sAZzg8a/31+npds+HaNDTcojir7dEcCWwnjk8PYnuBDW8FOwvG3axjEWBfcSUGXdb+Lk79dm8FLu
StBnHiBdG4oGdtFCL3NgwibnCGZAV9rs6f5mxqtaP4DZkgKOvyefBP5nw2REIFFyoQANxxacz90s
amCdM0J/LLnLquGS2KZ3wcYXIBsavhng1nbanhk1GBJDOkAIEtkjeKvypyweOYIkPq4Cfx0YvhWm
dkecyKRGy2IVDUJiuhUm0/9iVLhOXVeTYoc+4w9kXtPNChgApEq513DDf47qQOdmEKfY2cWP2KJM
ESPp5sMSqx6eXCtCzt+8hYCbLzoihlWb7RygIYOIvYz2nq5gKza589GErpaMDF5mQM0lY9LgNzQu
1msSKWbzGnU4NCFNyjINJe/QbWVe2EnJidL6GWX7rlRjXIyp8TEMvOkpvvgNwDlv8IWSC2lknwyO
aXiimFdJXE3T8afJOY+pJGihFAC4THGHxmEd1+COJUbc/n2Q3C0CaJACFFTJ3Pz0EN81V2IfTUnY
kLB25fhY1Tohy8tjZMdz2FQX3lg5NfRjCfzS+f6lz7S8TAqfDtgbgzqZjgeXmBZM9USKO+hrDAKI
7LZu7hslQw4sa0RDmQqbbCkzRQngVfBoNKop/4248iUqhd0XE0r3/LfkmAZzsxN145Tfb5lVkmOo
Eg2koAO/s1a8fhFlOyRRLFF95rCwI+18Nx6Dc5gdGwLyRsaS+KViQToo1tJWsB6/FAkJF7/e815n
62sASZMbuFq/z4jocdEn0tP5+/g0+ShXlJFFa3EnIPGfiyVCuQ8KP7/nZd7gMVk7aOnmPZTN0ls1
Ph8R6g5jESEBdQjjbc2uLb0Q2GpQSGVEpgEq9hjYtKFX3LvzpEyrYIhsHajggnlVVUFmx3hu8Y4S
tfJ7AYNb+vV70th/rBL9JcKh8GjJ80C+nBWDDVxk5qzelu3QR6nxGgw+mNG6DS8uCpnYodFv7E62
VfmYPnkSHMQ1NIaisjDW9z+B4YjUTQn+NDzW+lxdVj5LLq/mgu11fqeMJETOAIDeGTfB6n9S/4ny
sGwyb4yjreVavq0R8BtJpsGug1mLVq/NdRRc72bgAuy++jd2e2pCDaHINAJyRQXZ3R2qZ57ruBkZ
aUBTeI3XDGq4DG7yj9kasIRvrc3YvqtVDFgtIUTlCLdDkZqmGGJJ2eobRYv6H7BOEmF3tijwogx3
bpBRf9jmkK2ltKADNZtmAcVT8yt/PrCnuCebKLEZZMF705ICQLfpN2NQqrQOqpas4FEasWCACLCX
bmx2EpqrPcu3H+EzYAcu9lQJNm6izWltoI1agj8X04CT9Z6S4i4yNYQrWrJjRT0udtp50r5vKdNa
gnrooI3T3VHGkGofOTqqIJmWSNcpo0+7R6bsRP8/36iuYc3TFVsTL/7V4CXaWCb/EpTgsZE4sdez
6Qe9oJizReL/uUg2vC9Dt+2/UEhnRQcKFdjFkKL4O/YW8l8H9sbP/rIjaRVQ+Htr8JXzy05YYQSW
poImqpkXAZlTNBRJemwRjkTX3VxNBeGYsP004jTaQrnyeLt8H90x7dDOuMfFfCXFfPG+sXRi9hMq
oP3YnB5O79JwcIpdsv7KgoC5Z2jM6sQu0R7ldCwHJDuUxgry/Ecmo+Z+MDxybpat30MPpE6bRgXD
kLyv9B4AVc2RMz5gbt7uZdUXyKWUlnVDBqJW2OTWwNn3H+y8CBi6+WI+RVu9zif3TaX5Og11MO9m
ycoYHqIXfWUi0E+DMYu2a+3EDXdgCA61A0tSp8UhzLYzrjyloNZyHCFxbJFlL67mslAWEa3f3dsq
nf0yD+ddogbuVZxggrQmTmQYrhEjt+JE+TMWAR9neYWvBthEhKxywBE7aVOJoWrrN/iyXg0rMqO6
lMgzFPYqfzvNjQVrKdOI//gbJMbhsw7s5R4j9Iha7C9knGyFQZVe1+ALeV5QY7tAc1DbZ8aF3Ocx
a2cKySv2C7iT4s8zjWRWG0Nu1RS9HlSV5jfqOTwGouvRwzP3FmSBlE9YsHTf69+ElcAIWon14brW
rMGQclKMOebRUCiwiCMirSiNeplTvghsOQoRBn0Oumf/VZjMdVOp/6xnZSFMDXP/lnoT/bUryG1X
SBpLwlHilR30P54YNtUPEpseB0q1qE75q88zSxXb61OYNP3MdXLYUA+Zy7VkvjJHwcAjhindZXmh
XNL98dbdjlual8udrkLa/fOk5nsMsUAPT4FH38HY3YHiJWrpk3f/672ZOGKFES9iL9bZ7Km0K/GX
aPLU+YlggjgG40+aJMPCcBdfI/KD0HYzacf/Xdfc8qIh1VQVm31uQrVGW94ZN575/oLe2soAUv6O
JhRyGzHYtT/aEIF69ERDJwWhi/gWLNnIfJnoMEc0FoEZSjtExLemVrUT8+Jvl9db6WZNqF7SQNMe
rpbnAI7yNobaSoMYmNC8hFOwHMG0Wjbx5NUQz9j0h9ZyjwTuNnYpi4RHxm4HqBmccRjaV+HOjt+9
xueWYAWMcwxB1TOmmbiI3r3MRbbDCZNwP1v6sivuKo/Hl+jAsCD9KOwUHFh3vVY0sd+4fv2gt4SH
n7EmxO0pLNzPqaQvsRWe125SwKQilsif9crJx07L6nk5fMkDZ0XjeUIMjDvdgJaviC6a91IjUAux
AWW2iMFPWtYz32UdrfwsNYsrgTI5ER3uaFt39kIxBBumdIGYK8VQsIYdXQ9jZsankytYeET1Zb1x
r2zhm8cwqbAXWS+L+p5FNNv56IIVraQTYYm3oNgtAah+Dlb0/aLiRI39APBIIt6dgWD8tydFu/2E
xIyqGe7FNeAO8oGsZgBvjifinsUw/gSr2hth8hA7ovON8nUxLYjK2bdizg79IWVxhr0QTTO7j1Ny
XlmVFE4Z+7G/CyHXrQD1OkWdGZ2fJeMO08+vuDOFRgeaqKbRO8fMsJ0ywO7lIo1ZRkRU/ut20sju
9k7K6MzuFPtB/hjwGBTyidh/tyHCAktJY5jqq3yssWsPLrAraADb3y10DZ4sqnlxLCs/BiY4eBa6
BHOqQ6SckGIfPtTwGEm/SBFMykrWkt1I1YHOnaltrWqFGx3Ktr3i8jN0wzpfy0CKt3RpP+Z/RlKw
kSZEou2xFfEqMG/0cfuSLnKY0YV+XW50AoBag3Pg9ZJFnTreVU7WjcjpIEke3zbV4mI/2n6RXx0w
QJQuW19eZE/hfdQWWZSVEdou8UEEAbi58udwFL5uemsvqdK7AwreZZB29LsLjIFbQfqaFTRUj/Yo
LUnMHlMWajNkTNYqnogKP+xICUWiQtnMTMZJjsUAsvkuVR9ZjDyeI6k1bRZcLhkHObUDrYGe5ndy
5GkLXaN7hlMufL1eCZ4nFyur7RlmEKPyzpeN4tcbjyaN8SU4uZ0WLDYRocjknHJHfA5zCbmGWF28
5oHRTrDQKuxnJt0xRDDKluTtNKGwQUSAQJrU5N07Ybzfc2lz4VVPnIn8GVN+11AVlFnuVQsvcIxp
h0BQHGG1bs5E2gQWJtZ4GG9jwlMGlWROzVOed+5CiyYp4+A4KuGHs+5CFKjnUjYdHuQiX8PDWkVT
1AfnxKVOidsl2TllA+tmPKlJeN2xZC3GpmxMKjSYlzfY2ONMfNYhB3xe044DieuRsBKAlOVBwqur
2PeGuCilZPqOTsp+LFB8ME9SvFKs8xDxZowdaD3Ds/tRnzWGz4omL1M7iRNLrFqsxwsxeu72/Uwp
ZaS0BpzYXbtCoeDRlELqyOroU8QCom/hyrAmQCU17OWJ9LnOakS6l/Q1XAAbJdm7Lm8z46v77sQM
wpwREcgKquk/J0Zi3NiEpYTp75shDkacMMP7QyCmq+BVjpvqtgNLPqUuMv4WgEfZ4iLTSY2PPHpJ
NkT9xBAdZmmb/kAM+YVAQZuwFLk5Hd0yQZohYMFGKTAH/2RLBfiqYdZLTkH2S+50IMQV+83pAXky
Zdl4uf4zvLUjjFDARD2hi5nVLGpbt5XR1jg0inB2tn0DGRWXOhuVGB4kThKbI1+s8YA0CviCab0f
CA2+l/CB9I/N+gcFntNRbpy4df1z3zWt2aQV0SdPlhfkXvrxnwZOfvOe/3evBrhNYIAfFE1IOYKB
hCmxq6XmAClTMsps0ffNL6NZBlUOYhvQhq2TdLpfOmVkIiRENbtOGA3rSZAGmCkT4VvZ6aFYroOM
rxHqRbuRrZb/PD+VGU1j9Lu96mwKWcksGnRIHPPx0uKHu5DlFwXlRZ2aa5cfZxhFJo4AllDQgJ0h
Re5g75mnaWhjQ3T7LBmCLTpZm29xNGnIxmibNBR/H7iypqboyqbp5+mQzOpvZrdZjNAfQfrefh9+
y01IC6zzp8YK30MTBku6bREZw+VMReZkuMzqCHURkO2+2H7VeJ/5KGA+VKSGTXNFiPFse7St2FI3
oo7sr1PI3SACoZSV/saDWb/snUMRxb6twrR9xFIcIuudgi1MsORxzLKolkeKTU+s7Ox1i/GwPWng
ZB6ix/gmCQ7sk2C0bW91y+tfGus67sSxKDFuQIubFr7SO3wPEi/T9+CB5yJETggLPS3fceFJi7o6
mwLaIplHWGnegnhIGPb9kGbulqfdy/BHMsuM63lN7wWXz4zjG4vTlFfEXxbBQCUZdF3jTOCS9I9X
Rdm0iM7zpFGoqznuKiWBwpzpWlV2v9Y4n8TJe4q1oTRa4hP7pcdobjgmbDvk527uPcOn5qgRuLDR
RtQ5e1vL1F+likBV+igutpegugZOuXMagVVD1kPH8SUZ7B+9DEzcz+sypkyd8fVKabwhQxpnBeCS
L54zx8BvUhK0UoUG9KddlQ8hqpBN6sjc0qUVZfDoaToygXybBih6hon9AZivOsFAryD6H78RjIDH
oB/P+aD052tF31ebqKTOCj6AABKaBRE9gz7YKZ958Pi8vvq0aCQPsldznVj7eElyrnQEhZ3oyxie
cP53JiQKCvszEygNCCiCiDrDx9XrwejmDuJEXzCMrdL1eIFtzKw+Niw07Hz/5y+T64fWoWc6vH/9
600sfKxw47k1iwvGvRyfBP9v7uPDNRDILM8q8yHu/rdD6KwoUTlX0FhEjP+55Az+4Wtq7+LkU2K3
/QVFjtrZdokYt7l1PLtTRHSbBv4ENZNSQV84PWluDMW1zThJYyO3MtG7RvXpBOwIPAFK9hzb4N5W
3a31PyYw+nstPEcHF6aHMvdYfom2qsO0136u0YF6hzwE7ke2RLxhC70mqJbrBGY5jdH/cuHyt/zv
fPyogkmONx5VzjPzuVJpxG04u1qxMcyJwuW42oB3fmb/3q1xBVCz7f7pwqHn3zYF/dI1pbwRFmyU
/GqXRhTr+o7gbMwhEuHggF+T/kAvLwdb5Ef+ec1GppiLuEW18G6haVKWgTBvvvBWe3krkT68iWyx
fi15vnuoeuvWaX1WMHip9NC1yRkUhqWMwgUzhnJW8vSfeBJEut17KUCBs1yeZtucaxnsAQ+j7x6t
oHyTY3o9RdWd4Roz4VWTDAb+zdXZUDS4eJ+ORg7GmNSRZLcrdz1wbDn4Yp8wss0Tv6FQwM9lQ7r5
fVgSB2DbXcgtTQHs209bFRPvhlRk8lb4VIHPMSa3hEwjW/M3JvXwZvo99kbqyEQ7xd3t/7FT6c3B
g0ewLBW+9C79heBp17XimcP3X7DHV9n1qJ+7Xro8TwyFkgX+RKJEaL+ZI1aZXzkOxc5KKY6VKxZ3
ZGPeWqYlkkEBeidmpcXHGJAMYvchmlDyI1JLzcgUJFn6hFd+R2HdSppsziKo6foFTj3fkskyE92g
56ChgXVAAvrK3akq1JKxFlJToE3fh/3CgRO1ihrYYE9/W8od+VZ3lG5xoUkDP+7/ELjb6DIeoQgO
fTDKnP5W5fxIkTRNyKwk
`protect end_protected
