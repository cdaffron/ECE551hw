`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MbQmMUpdggsnpfF4Z7OtGUnm3ZkqnfpZFLVRZL8onSbmaUSy6A+sWVi2Xbj6/C5OpM/w6jJ6z7DQ
Rt9lMyTeBw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oY+sJGzyOyyczoyALWVEhEmUaHEb3YlbxW+84YQSal4aB0Q6BVLIH5y1x0O6TBw779v0rpoQ6Pst
ivtYSOVzD2emegOAmNNGZINqhcj2FXaS6+y0566KRiGEKKzUILSllR+P2WbX4Q8igKUYO7SA1h8e
aGpljiC7HV6222Yxi48=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sIBjnSNnJCUvzcmwo5fMUZc3irEqzyCRlf2qcpU4u4UFPko8/4fbuPFPReJGioM3/dezpSCOUFlY
R0qJ+9aIsenU3i5E+3NhFmaocc7LlCK7T8efOqTxQNJmrwOk2hTrTy7KSXE5E0I/3Iyp0I8guIYs
/AJKoKF4tnVubr3WlalGfWRuJFi1pEYbebu28M6wuqADiNvtNKwALNQ5QV31tLmZPj3Oq7TBd5zT
UQRtCOdJJQxHWLlHxfOJ3K4GtF47w2OKsQRRwz7GfBi7dT6yfAOpcpTdqD8nsNAwS4cEP3o/lkm1
a47r/8xC4q2fviR1GGed8TwIteqdea58XyXkSg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YfI0LM06mRsnNfA4qyTxMAfI1MQ/uK1Jim7JhF6MGXDYgebUlq77PsCDoPznxboF2xp4DV6YCppV
gqo0CQP0a6zV9ZXS3ur+fqtmFhk5NkLRkBu7X2ILSrYUOb+0BVCi+hljXtTT9CVNnT/nsI6RAgi0
myo94WpxucQ1/bB65ZM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F8OQigkBRu1Ccs6lenUfeG2qddqP/GnscnladyQlQkXXN08uZuQErcAUKHi127xLkLHH/B7HRC0x
Z1wxsCyeDu72OlU19hqjQjkoOx9r68Aspk1sZJCGyiJ3z9ld45yaIanAE60LLoXMRMEDb1kG1tur
h0cdtX9rOYcEWNkmz0FTisYPstB/2E+FI2L9h/siaCGGUx7RLhvUNZeEexGZUyL0lW6f96fLscOM
NAs3LZPXa5rHAFe6DMBe7iNb8KctQOUHTuj0dhsyAmXwgJoO86af6An76pTf90VX+WNZk4giTPLO
qbZjjCdGdS6W81RImIGjYw9hvOE9VDjwyweVKw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 156848)
`protect data_block
6Fz42YoAwiK7T8Rv4r6W5r0DNHoUJsPU6NsftouZLIZSXFzpTDAL+D/YrbeSWJjust95NgyPxC5R
pDAa8OZpIeCWa2HLMr59+Hl7etL5oPhmvqoot88fnUXN9NWKqoquCrL7/srJyniXsZuCo69pjUAa
CdS7sDphgaG8owS2WS9XjsWD6ONEkvFm2Z8Dm4Fpz1tdW6fo2wtT0vO2McVjpggcA5pJnEDqQtDb
ZE95GVcjIlBF4Ag6gtSYiyxHpJdX8HyUhJJ1VDChUDqDpjlejJHUUCVszRW+I2UlQxuY3c8Pzc6c
Z5dokyIIMuR4FKFZy/s9Jp0R6tDU//9i+X7m7mZ8Eov8KIWPd0i6QMlYEmINTwo1vVm8SNYqZzcN
kfgI6ysphc9WOPPBJkecU+zcuAwBDe+QNVbsCFsiYRCXzsp5Xm9KxAi+OWD5CPdohMdXY9zr4u8X
+6Bwf7n+7OSUBMw/YZHNZG9DH/oeQBrHmtDv9IWuKswvACMaRyj2MCMIxXd/JhElJ57+es5NNwgh
krLTEI9WmKKuNZXXgDi924proSAo9fdzXohRjMZiT9RAtoeuAFfZW8uGUt2fKmpUTkRWhcVz1UD5
GV1sSdNrJuhT+gbBJdJ+DIKB2wo9/U0Lp6MuvdWi/uWoI2xRts05P4ukhaYm/WThR5jZmPKhzQp0
gfEe9vJ4aGVz+ROHRgZSAOiXIdxim+CZ1xfu3EAFXBE20+5m74fHC3dtFTWj+MjjMgX2PDE63sGH
4tOXSI5kUGGObi7JlUSRlULjabCxerbx2a9fWsViKo7j+VNM+s9e5y5XyTOOP/6QtZ5M9Hua8HtA
qCxqGre4VHEPhN2ynlaOE+LHQEbXvNQVHUMzfZTn+T5sxem4Nmmguy2/DzoJnwZ8/3KSPLtSJ+SS
yHTuM1hvoToTeNtUThvZFuCOaZCWC8hEG8WvO6chmaty/hqD5hlsy5Jq7qK1gEoiIgCRsSo2hmFC
ANryRzLEqwhdcWbgGUhHvej6ZvYL2l7pipRzLOQOMhXRBAkk4rOQzMv0fcFe7iQVtptWOv62GqBM
Kqir+94N3hFgWCHfZ+ZXjg0U2tmcSpOtRap0FN4ipq/f5m5rqe/BV3ZA0HxZRmnewITgRPNs51ni
WjxASsswmV7tRp5nbU6A+9A9BVJXbOYC/kAExWnRhM2tix6z30NrrhqxoVe3WKozNLzjVdVMnTMY
o4vLQ7rd8EeXJRIF4xXembHy+zudwthwClSr3cOz/4SddCrtq3pVPzJRRqsWCW2doGBIUGaGo1Mm
s4hsgjfeU4J4P7/w0vF8QG8apdKD1k6+glL5FW3NYAhuoLE8qiIfpTqMeCzZ+YV3lIr1omTVxxHx
de+Gj2lwZN3hTnzcDrnqeSEYj7990AJRun6CQn/OWI5xBQbS/ikuLHwrs1Riw+dQNbXTmpAwykZD
I1DDz7mTCX4ozrZFjiE5oYdzytXmkt0Swiru3vZ5xviN4gf1k2KqnImomUYayxekbT39clmOokVg
R2wXXUQ/IFJAbU3WNi7hF3PzylK6nw+dAhPMBkFgy+Md2cJs6tpzjDI6q8BSvPUtr5IHlI0EUd3A
5HWoKK3W5Raq0uFG88faFiQaI8MRH14c9JLYwCa8xMYNgGFeJIfPKZAuSHtj3e/xjFLiRM7sbzi+
FEYXZB/CoxOK/m9DdRjzGqV6mejvUyoJpJHsgQBSAqJ9WWBwVVFhtCZExaYdO+ycApGG7Q2L/Hox
BG5ueFJ2C9aKN5W+3b3mPDm+LhQTLFo8KGC9jSWELQhL1I9M/ciWoE9vA8GDybJ/XelI+b9nyLyM
7TLM4iIGgX4LdgzhBXpUlIJdLnvloNVGxoJ7rPnHWC1Id/WWRx0rB34klESUePepgt39qVAwwywS
AmPmKw9L43C8Hr/jEQ+S8DI1KHI9GmMmvOPsk81KZ3rTQVR02bdFOM/OtKf4eOly0IHA2fpS7QjX
NGawxl1K+cGU2mdS3Zo7tun0RseSTQ50jrVZNU640cS0plSWJmLTP2DPDNk4OxIAVkibREYQDhI8
vUxHqhk9SrscXaMsrizzeF1K1daXBKforhAZcjB1CBPoIOK1/6EdBG/CmCQugd1mvFxaom7zjyLL
fHKXaGbjd9s5QTIO9jgeFtB9LrNJtjue6FPcEoCv7n4imwlzXT7lkEvUf1/b7i9svWfr4mFVbcNe
vnTndZX3yOFHooriKcLB1k/ew9qt1P+XowLLUwiQF3iKirVU948KnaueKULQUlQpHuzxIxDpH3PH
BeQZzniSPBnqiuU8zp0BvQdvuaKLVmUj9L1qCu+OqrN1shqrG4pwQWbhdbQXy4iHGZbW4i+O8So8
C1mG6LjkheF3r0aITgZIFA0TyYhFJbNOCoCWfgD1pJKeif1SaNRcAbmmTmwydhi19RCHCuM/caGP
54EO1eSVetfzjidcQCDJ1l68pLTzY8+LwO9Ehwvc7mCKieu1ldL8MoENJT3BRYBiirMpFrvOeBMW
bP3yfk1Wmzt3hZdY/Zb+wpLa09NXG0j8u7d6df+pVsH7UdLPUxKvjkoN6PIRGErfV+m1Z3T/C3PA
0BONWeC+pFSUD3jwe0NXrmSelEPubCK1rTfPW8mgeFOejZbj9r7f/WKhbeq53EzW2SWsTaBlEwJv
49vMRaFBUreOiWU4QAYkMm8bbVueuHySVkyl7+ObXUrigTuA6Bp/Bcuc9DNLfz7nKy/NDAAjQO3K
ESlz5Xh08uZpHEeHCxqttBf1EJrMkcyU1BRC24TMz5Elk4t5YtKx1FLA20WDhe+czHBPYkEcKvGx
ohEMUFFVB7xymDrE8PygmhAVuYSBbTypp9KvdrdJj1OkSPyfJTRyQJqgBQFU3L+LAXUzjNR7Zioe
L0577il0OQW//W1RBRXbBBzlT0F3l7X0DzJ5SkQ5CIveMkTzOmrULkSv/co3fKLfj6MMTNrgSis5
/jw2cHE85TsBHTLB1j5G1q63pghhzkGMt/mvXoNQNyXRN1S4eqZErXw4gOIsLqwuJbfDKuFo5e0e
PSahPKP5gQtjVbR5NipVIrXhuA4/gmJFRQKgKYK5oZ/+/LfVnbEG1AVtzRkOCG8io/sS/aupcR97
0TnrdSmToPNVgnRCmgloLwjdpmKJQy4V6plVuLi335YOSqyt6UNYwaIpy5Rla6VDj0MkrVlTR3ek
a67oKhDJ1s4lJZ946AyTCaXpBYcGKEeo3MQ14ot2PZ+RKjPwTiHz5bRbvQnETvO8ZSvL600h1UWw
5FtGALzSNHiypc+TfYTfqtS0he2cX3WYUgQBw1bb0N0quZtfMK/5qINAGUuS/c4N7tfP8+5XHcIm
d4CfCKeuY412rlbVxW3ft6Nc+L6bwj0Pavr29T2WSDlg+tQQvW8MVoSh21XsfkztYMJGTpiTQaho
ZuWA7ncWcyCpA0+JNBu2xfzYbIGdAjkrAKVR1ufgqMJs4OX4oUmJwy9KLcj3mAKkPJOD2lcd6HeA
oleYo+AsDsMS+oYHiXzb2r55ixA6uNx7kTaPmivtJsbml6MUxeyZco6dVF77g/3Wq3JIclc0SQon
VsgRgn1CzLAobG2AbQysD5qIwXHtlViWAYdnQhu2MAB2PZlM+m+hTuDpf8y9FYLbqvMhQumXxCGv
wbPYfhHUeW7OQ9osG0Wele6c6OdYZ1PWN3I/zBSA8HkXwvLTE4MosUvrw0px8TINSCOEiFA4Fi5X
HHMRyH+Jiumzp0J0OTEOC8Wc4EupArn8V97Gb7NCZfCFiKtPU3LLd6R0EQ6ja1vJGZwXJpcOy5GT
a9osbZpF6KP4kHmPYPBNvRQaMTUJfteSUKFb47CV733eAWT+XNP10IhfZtc/42OSqdtaYywN7l4J
yNWrBIh5O7TQJOq0L8AGX9nD4F/QxgXuYOmnE0i6Y1u7yGPlTL1F6VZwMYzlL68yjram0n3oCkSY
NScoLL6xT8j6CMoPxS/LIx/DDm66zHIzvJkbUA/hIj10iA4NspDdMy2uCgU0eNotn5zKWql44XBJ
RYI/V4Y7V+PyH6Qj6knWrtc4URgx4uw6PZd2gk30EhUmPJ1qmbBLqRwcGoC6DdSzDTsezN3HjWq1
2aYrZ9D0mpNAVHMNsdoikSsU05S8JBMVsagwSf8Yvj+IH9hIwQ4VxTjA5/yA5iePz2mDhsAkY79z
591wvc2ponAw3HOocuymKXRsrPwFkZg/+AUdbPz7x1nh6Zi6i+lxrhzcUdVk/iVe4X4qG6Um92yx
jIyQnFwgEZgSX8MMYzqAYy71Kv/o8T4hWaluIDSCCcrsF/HKbc67MS9eEQSZw6m7+tME8iao6ifA
/zO+FJPhG66iGPNW41GSyBKXPzlZWQFxcX51hJDDAY+lTzPknVC0qrfBH7m40lyDYuQEcNxLBuum
Tt3QenC3nw/uZSiA+AjtKsBQMLK5mWowwtSdvjpsQzb6hMtPfdid45faS6YYF3MfeXYWiy8pX49g
1EnyvbLbI5gPNDalDbhIW16Cv2bumRHdmV4UG5Uq7ZU1GYULeu2zeMCg8fKgQWN5ciWcJUEA1Csd
LlULuo+Gfc5bVfI85nfeUZBWzqUSpWu5E+KPKL9SW7YIwUOSd8iTZQlYpX71d0zUMouvwzxB6O4U
ZCycdzN0aulk0PlPkYcYE2eaMAW2sjR7rU01i81ollVoLSF8g2nr43HdwbxxfkWTNfgBSailZCAV
5JynLPmU4V0ZsiSMmxzcRGAlHYHG7rL1XgYIFPoX2WslkGTl0xEMfARo/7QpiPKh6eXuQcb7qH7N
6udZxGLd0dVaTg3zhqL8NFQ1MS2F9ddAaGgAT1+7ZSx3q7TsVJYbTltfBe35h0s/zL4QMdIx6gEu
Um1ntVqqahkiEDHWDLUzbITGmTc7rQsxTfyX3JRirwRNVfaBdriak+Jaoj/siDBUdC3K2GvZmUI3
dd02OCY97pExJnB7lcxoCKka/Y4HIfL+Pea/mSE/1BpEN7yYk+H3krSmhiSTqBFXOr+D+3q0Op3N
raijXUCOa9VQeyNSE4QRcXzNhNLqMsxIERyHXI+YQobCs/cmaEcd/e5Qy94byWQ568gynBOHrMKL
PUNKUilBM3ubfvP/L3wUBxRqNpnvQebOHxZqdmovAen83lYXeGCOUkRWgpiNyuZVwyuV0NYZPs8v
zRU8Eprwx5wlOY8s0Gu630T6nMJ3tUw8LJrH7NnSw5QT5mnTzlwIt+VxfynZjVSwFW/wKfIvYUI7
RLagT5MKd6w3iPzA/dySRLRjopInjrEc9KhVAtfa1Acvv/2MZLwJe+3HInduPR7xsWNk+O2hd7Wh
hThci+uheoBcBBpGqHaiWnR9fKGZF6YZXt3s7xYJK6MzIT/6HdZbnG+isyINaf0OxQVGusSwatL6
7edpYiInMXXVVdbrLzMrKn+loU8/cIH+C0CQeVE5QJple8KabxT/Rg/XPI2AoHREQNCUI95f8zRt
nsrZ2yTQxKZs/uAgZv4TPxFxncUjZxmuvqUrqF5ohxsmZQmLuYF7xzWRi8RT4+cJsnmc5FY//lKR
XuUxcyXzRkzKIvHmJDcSX6JFxJBGCWSxnJqBKXvE9sRN3fgJgEoakIeyJB8JtSQeNXKf5kyKq7oH
ZKaZMtUEiPPkfTa5bj4KqOJTNCWIDLIMg63LmmHsGFFCPl8PrzE27nhH7Ysaz9BJL7owcNGxZRFS
Cb7mmY0dZka2YhPpjFST0QzzcJI2arH838eUL/lFZL5oEAsMaCr7sXmbieDbDPBzksmTpMnsYZPj
i0vVFubi8Zh4gATpiHUb/QXhq9c8joXhjHoyXOt2P1k2ieSKSfufrmNeDV/FiU5s0gzYRmmKNLEg
YKccd7IzSm5Xdq25Wh1ZR4Ag8BmJ1zxgh2OrtWw6MPSndyuliw9AB+pWNKpuyy7c4x60zTrI524j
wVSP91Yg9EpzSMwMCNndALApUH7ZBfuj/FjOjunBtbODGRU+uZhInwm8tKCRHORH0FjGzOGFtrsn
lfPWG+o6TFaqkuLb6zgBxQvQCHDC9t3QX2l5XM8Q2gidOqbgCptGFjMhLJI/ASBCngiwNTBIVEfb
ZF6rwUhWqc+tqBYYFLfZIo1tvrxD2NxXJAuNWktDzX1lI3ZXBbPcseb8xCbGrT8bYS3pcXVKFjNq
UaZsIDh1Q+f8bI+hXEWgj3LM5+Mr7K/lFgYw0FgoG7g/4xDPDnWSTKPjFNv+boUxm7YSz6aBMdCw
I1SMHVZHMnaR0xJqR4RwkHuza9Ds5qds/mipyEijtvbmynz/cQ65r2/r5cz7f/wIz9ABRsuZ/RFT
XVNpbMv1+D28wgqNFEviWpUoJcqYrgN7vjU24et6xmGosCulZastEV5SfbQ7rcH5RAm3arxV6Ulf
mpRHkMZ7e/+Q6+vMOn/behWc6y0017/7jTjq/mm4lWzZoXHxGp0n3oRoLGzSEn90aauhD8TIYHhj
NuQ1X4iaGE1uCWlop4sXfxV/oMmhS6saaMDZNSa17FeCVxZoYadr5kjRSbE2O7vMQ5AxuwkjwIy1
dvkVn7fwyO/FHdqMIcytibJta4PAXlSTsb7OnIXDe+Q5gKpnUQjviGtuhwXR4w2FKRvaQo0caHkZ
RQllmHWlgRD+SVJLKvhC2cONdSlManXhgrX4cNLqioe90cYcdL94YnQQgvde0Bc33u/h7XhEy/0C
idEsy3qBz805ZIdsTJEUTre5jPtlAVBpyrxp5vVozSz1/J5iqUz4RN+wrZMRXrwCW78UXKoe1jhw
B2wjcAXv9DMD6HbXL4M8Mlru2Xevu8lI/Y9ZEdKb2JAsHsunnJSIUAwCLdOky2SLLchfQwy+KjeC
yk0TUBOi2cDjdP0RULvbgdLRAJhSgrNxJIcZWeY8+EXk4cyla3aUEpgKYGxR6tDpD/MMmVE+I55M
WWwBy+G1AziZsQYG3/4pAN1kHHC4zOKRKMqRr4G3AM3QoU0RmN8iXkBO3VYfTA/zPNWA+p3kmwNv
8vmjf4qU92in+6kgOjjahUqwYR/SS+qn/vygHXHlUhfwqceCVQG7XZ5HSPKmsJzu6H0lhI8unGiv
8UbW0kTBuk2A6BJ64HIauPQVGrBY+TX3nVvr6MyuRjvGFyz4c8/tLgbeMN/7xtHM/SfOy69j5hHp
pZot4jFANWUgAT7IDAvXvFYhCzXuxJbM3leFIvDZjp/PIw9uwchoKh8ccWZUmg1PNY7k4qzK92vI
RA8onJjH4fKdPfdWp5IKtldwXs6urfenv1fBpqFwcssJXh5qQjmm0KZ5eV8ei65PYGZFE3R+AKmi
DOWUCIpGN8mNExOoK6bOe8vGAliaaV6rLCYV5KU6+qIkBCu/b4VAC4oTy5t6J7INnRBJS81Vnw7x
2EKGadRg7i50yBP9AQBB9XbYiMdiAGTQWWhI925mLmw4tsgBFKtlgQbLolRZC30zi8AVKZCS2dI5
RwbWb5yy/23gAYS63frTr4ujFDiP3ujlWfc7ovSwnBRwZq2PsCG52cMuFi9MIP8PfvNWGWB9GEZx
t7PimRZxHctHfOBCzyRlD6yBPJEZppDNxkfSdTNlXX/Xqla1iGKZmeVxkjf/iqEAuCVkPnmajjdD
wVSOgWB6t6+j5HpFOdsp8UHSLFx8A35j86Qr91/S2JDZ1yLOb7xmpozNYukfjYa3Zr+I1XvBsIt+
tNvxc1TG+M4AWENFjM9WYELiRroQ0Cbnfr3DNN5SWN1l4kOLBU7B8LdTXRznoLIbGyvIR/48YQgS
bwtOVfREtxnuAd94kD/5oCo2I16lNqMmQrU3xBGYPtPse2+9y8zQRM+c8o7lMyPy7oDRLscOtRnX
sg3fpQS/TNsbhrBnP9yi6hCBx3kvJDrRL/uvAIoUgTli6FGZr123/oY9oFPv0XgD7aOUJNcdvHZ1
Jb3N9/th4HQYb4ZDRzLklcxS+iXUckzTKLW+tZE54pMHhIh6F9iwjQjsjhWUoRjGJIwGp010V7b5
41hnXWLBsDvi4awFqY3gVuC2HPwOnzy3HLKLQvyTVJTjkQMSfQFwWLpmaG8/7AX841HPZ7AgUNn9
CuepaRDZWnLO3s9iDrzrYxSxyX+9sMfo2NjUai6olMN7DvgQ3gGz2alUAILk0ljR7gFHUfE2Kn7T
fGJ0jffiAKy4Adxgbuj1QUwAtCIs0tmFtOh+SqcNx6rXAdgN2LzWN9ZEOxZHRpgr8FVtJXOtUTr2
+67xU2lH6Ob3YdE+onF5+72xwJSJUkg4EeUP8fSs6Q/l1JrqY0vxY6dieBxX30XqVISFiSHLV6sI
oS/++BkNqwZhY9CD1aAO1v9HsNJBFVhGTwMZ2owxmPBvIMDOC5p4KOvWYmiuaPhYm59VRYDCkwvZ
kLDo1E5PGUHIwCDh54OZ4uR1QUoV6yCAF5Xhi4dbjq/rKr/79blHgkgUi0CrKGqlMgLITnkvYp1C
h+OFMk7NcDioWew1oZ3+v/WcEo9mpDls31bwB+NtKz5uIXx6+IfwtFcAo/aeqYnG8L8PY4kIO8QR
7auc7WeSeP+iWA8xrhdNZob5ASn26XYPngu6N1MDJ3P58IG+jxQKXCm1YE1843NWTeIdIcaNQFFg
kcRokMTFAmba5USiiDilt4ZYcR384srKATcZa9zFj2Wl3WwJAz5VXDVRhhJs1QqI9u6cUXooSOIm
JmJIhT5dg2jkE6GQDh78mC86vTMBRwGJ+OJD3T0oU69y2WWpMkkXHHxMzFuRQb4ogpnjQkPYHltU
9FJXlgwk5rfCUzh4C7by+jWnYhoIMu6jHX9QQsS5PdZEVmy3WOnFKqBv7Hqa7s4y1xXANCs573lW
6pyld2EHwCruNg9uNwGdVn/N7SAAoUtHBDSOdHcL2VgsmGGan+W6YYc46LU1ah9Qw2p58Ey3hqfb
yKVVZj+vtDS8AEV4vbesJAGUPQLlm0V9LcN1yvp2Xm3hGXpS1z2KrGrUU8t3/PFl6uuSI7xdGPgE
F40Gvg6O9Mo4y4ZZvni5ByqOgB1fjFxe+/QHoTbgDTW4HL12OfvgyfFt89K9PKFO2MLHtfZ0HTC9
LebjNtQ/svbCwV2l1e2/bGwSuh1DUrvPrg+R7ZDEQz4fjErpnWwQp+TVsL/tklSSHaKGN2Vwmx/O
CubXXoNmALdZ4v7pC3k/asDxBz0Ti0DZl5c81b0EO0UvFyJtcmY0VApeGWDTMqIPjUc2TpJujxC4
etMiKzGznUtiCxXNX16NuNJloDALZsyAnzzHvsxmcbdGzFU+2ppE5ZzLk4c3WStpLLxPGjOU866g
0MKNfzVREN+xD7IXWAAK+rCiyuHUBgfxmKN4gQvzKf4+sdEuPMpJ0cKSjRvtLe9BEVL+1s48EP6d
5vOHEWHd1K9GKZinwyxTdTU3ZFskCxpmuSkpJV9U0I5ywR4iozktXKllWZbVH+OizGlGiVSFhokJ
zlvmPF5NEdVE2y73zKsbVCTQkj+BVN80LQroMlUioLUkdsW1yQ581WKmJz/B6HBdl9eyjK7pkt0X
tCzF1SWKnyCztt6iHzyMmztpatoC3MYHLBRSt24kUwckWzON/W96oPrkxCQM1dsN5dbJzDqs7wqc
UOLDTLUW0YiMwyN0szg6UEQvLAWf/jHdX2/7YBv9ug9rYEY5f04zdsLpr95vWzLsOh+vs0L0wFOy
U1i1Rox+0uLchKzkNeb+nnarncxHnkZTDupSHFT3Fzgy+5KcEcP5BHTh/2AXZhgh4CneGQciYo6j
t3K+VBQpFgHK4EcepaeAJKvgm4bAykMTVA8Egn6P/DvlMF7YiMLerzEJL/shiabbpGQuufnYrY8u
W5QpYiAgzGng4d24wRo7b2Xi0jCwNajAtDOueZ2frrZql4B1UhhhEa0msZzdRHHRycFqp4XMoLNS
pDL4CgUe6iE1ZTI5hyWT1CLjQ+JLVNuFyRZzC359qLJiaimx6qZIVlvP309TK9T5E0P2VPxvdUnT
bHWVXWXuNV98knpT2KChE9QVbNwvKVYTtz2fJmNJWHuHrXtAFer4aP4U4QhHM1p/ii8R+jubMEyE
iZMkuBKnoYP1aeYEDak1gQP5zb+v/2xWYVdRxhiFHyBUqzUHa8DAbDj1iEEmCwaWB1cXPZS5ORyg
RYjW2b0z+nKieTdGfynGZ7NxtKLSJT4eWbwj2EOUtZo7XWlDitIrABw3LW19q/JkxWyJFPYSD09L
fdqWx65D6nsLXeIwKdnjkkpxEFQbL7ozJtR08VuredY0/he5KEw2g/PpqqK+NusLe8xIx2icsvXq
2Oq2IgXfeRcohZdzfOEmeAgtr3pQ1j6jD8BIUgyFLOJ2pD3jyNTzvK6QGJqqAF76oMw3glCqDqf6
I2dt18ZIroHo81DhVruNTOz/VZnQp8XpE3LU/RGMoOdk2kWfZs/Y12uXoSQHc9hP1OJ/SXETT9w8
VKMDnbnVcB9U329hbXIBSg1AptghGo2aso0atpSVvPtInayBnBG0F/t/07a6XZRxdZ8zXj8iXAUZ
dnr+Qk2dVQAv1p3CezC2kK/nHbydtKUoQ0US6KRM8my2ADG9bG2WKJZGZoRF3pE5BLPvC43PAa+E
Wz4xzotfi4w9UZcBAO5ajcfNlE6Ge1o60mK+qoyewqmGYnlTMPPgj2fnYhvG8UMtCYGK6S/NmDLr
MkzvhSmgVCKIkYQePdAglsnjkWSwqy+Nap3rAWWpX64GrkBF71F2pNDsrLGwmgdb2HgFA+rSK5tB
/nmILPRFRMsjS8rpz2qy0dfZfsoO6wun7b/EQu/LlCxSt/jbHr5QVWmnif74i21OYVShThBxS+Ug
PIAuQZzVX8b1px0YXznLb+58vMawhMEFSkiDjuSOmMW8DgWxMilnrUyfaDDlH5U47fnWwn+BIeBr
jo0OP2zqiGwsHPHFsCksGbvXMJXFvpL02Mv67ojd7Fl3oq1hnhzscXJkeYbjNuVcSntN9ik1fGta
5qivcjCHQt355FfIBvCJqDgKKbcuCCZ9NeLevwvXzbvFiE4H4cy+miID1x/Z1pqClPHK5D0nINUt
oeBtR9NRj3TQnI96pO5isgZQbm7hgmsJ8kNDY6eUahxx1kpUtWqti+4V751KD0hsoEd+k/+CDtup
KM0h27CvHPeQy+G49Jluste75ZGqep+XZxgVtYp52VR1WhP20oVD4LTyn+DpmIC1KHIgGO9bfylb
A1XWYez7KwGk41W3urKCh0ZikffEJckKrGX738J7NEMAc9NyNL28ZZxolqxcxjlTga6UqYYwlaLY
A1Lz7bPnxDJfkcTGMhXSEpTgZWJAY2vc9HD9AMvcFQ0TuTanaOZQqU4EchJfnYXbu5utJfFMxItA
2Z/4Ia12YECQd7nb5cn2/XhXwGbwSqNdQWS19uBygnlf0AqpLCAH/UN8V7ssZ+/dj/bE1DvNHuYZ
WUbdS8mMhEnihPzL7LImRZJ6TIYsaIwIuVLJ69fiEmaQN0XkZXO1ZeX6c0QuISGIqkEd9QlfMWqq
Pt+gP3+xhpQ3u3XGBkIKgYt0Tb8ByrBuC/giRqtT3DruwDDr+6z6FM0OX8e1xBGLdKa6274T2qSm
UFb+pvPzyFir7Bld2dybAFJNA6KSz19S2izkmjfDZVenXvxDRhSKW7YA5UzsJR+wv48xS3/nWLZ8
FYR9ygOcRAZ+zaZiMKZdLTXfDFIt8c/RfgIQH73T5WLVXiN70x/YH//nqjfh2FodRFd3LU9O90rM
vB1vCGUjC1gQWXV+jY8nm/udNcYsYBaWkh8TSqZ4RJq3zrXfPGdH8SsIeDGbULnmYu/wdYayMfUK
GbFIBTqN1wk4pkZCFGOSxyR7NLJ7C54ClIYZ7AFSwzOtqQ4UfwMkhC1MRU3SI1jXOjHMktUntOMZ
zEXcjxmoocjv90dyUPAKDwUlDVdtXcgywOsSaRx0thPCje2upcHmDhtpbRYagslSRhZSdjmFTx7w
901UCTMg5/T+cAv3PiYbblLtgUHkkt2Js4w0k28YnGzi7vlq8EctIQ+eczB4oLUsZtIJFexgmpDP
PwySvmZUjN7CJLuwCUY9MgftO2jX8ssP6qnogJT8jxhrJ14Dq5Wzzxqc5NUBWjq66N52oa5AotYD
aryO++ntVbLr3TTOHq1585/BABkVj9I7CinyBGunuLxmaNLGrr3OfRNtFHa9T2VgRJlNMRZtD/5I
lt1JJd3lADEpnuYRRLRGECS6/8s/gyRx8PxVC5AqiAvak14wWKl7OWxzaTDcJydgx4voWsFu2PHr
rrG5P7dkT7fCDLDfiUdPDdW7Ku2s0X9iwngqkBGT6YbWLAABGj7OLtpHOoOzvmesvA2AcNq1dtel
Nh2IZ7F4762G8+41qN796a2c/FFUicAxjQRzKlz6Vl50I3sJDB9ycZ4Ck2lr3WFN21i682YRDi7N
X0j359qqX3Oe9tM7Wghgt7sbsJPjwfD3C+V6ZBLBWa/5Mcg/YPPxQ8qb5xifbt7wqS0Fm6Drw0ad
Gfl1Cgr1mRqgscxOTp2wW21Rxj3FdVYKNxPqxIiSaX+ndUVEkny00N4ueUGFy9EpVdjpqvgAqNGY
UnWD9d9RVuy3ogSN4n4K21lp8CtpKc/OrHbDgTGB/kvaZIoMU5i+oYRdct6dYMgrWn6s6egeB2HI
szd+EjDecRbM65Kw3JTjffrL59kKCLaVSqIDNF1YhGWMj6SGwtqXcDZzHWEQZWrvQAtCNORbeDmX
5V60zKiS/DBITfaYycX1Dt2DctABwaPJFeX4/vue+WVLI4UO33jmCOzEQSannbeYMgTmWwftrLjZ
jF6gsVeVeuTBA0+BPmri6rASKLNn8sEuYQrLis6nzlYWV7e+zWYSm7INV+0ohZBuIMbPPtg/WPM/
uIVtVY9bY6sz0zyllKwfrW4mJlKbDKe7EtYaMzvK1WOSQqwBsBW8XsMx/LhK7MfjcNxlTvOUEBM6
4EaVnTY7dI9F4/pIM2cciTGONGrPipgo0ppUvEHbSXyy50I4yKl+wjhW3dpQGiy1xnfpHpbjZmfm
ubhy7E/uALSIF0JHzWNIzMh9qEgimKg1DKSeEoXTea9d243RCB6RsVPM0noS593T+R+5viC+Ng0d
7r0Aadw6/HKKuTYF5TaeRCHkepr44JQlfiUS0Cv5biR8lLb4A0kfGJ8MRWeoxiYN7uoZ+k+FFv56
pYA5zwYfN7Ut9mX4TIfzc5qyN/M82HngveuU7kzNhczGZbYswscw4VunKc4fw3iAGl009yMhtVRq
6LwNEZYVAEDHfcdQCc91JRsF5m3BBEyw/PCs06oPy2bcrKqkYKve2gLaYmsv0K3q+/4ylVuawkKn
bz2MZFzYtTwgINoAiTU9qTBa6nYqVhWg/tKFjQlfBWFPAKqvDlW7Knox+KppCpNqwQTgiwJFm422
KpsXtf4MhafBG5law+lmBu2LAOmzA5h8g41YhwESf99pUAvQc2bdwWo+6kOw+vl9wQ440IHQM+xp
wqDsY3MGnmZCwyDa9iABDGzUQZQPxCy6FPeIx64UGO7DM0JhqAd1Y3HpVJhjCvEqemEfyGYAtglj
0gRs81xkvw6LlF8wyS3TwNk4MM3MAxZdzxQEMBQNYeOn5tYtYoKOHRmN+zTvOPWwQ+8ga+wxTvCA
AbbSj+3cgERAvkDj6/lb4v48Ps0ODY3bbt+3oI4Fu671Jn3/yDcGXSegcoQ2AK+s2DpymxWAJGKg
cwh8IXQrrbvdyJHuCLGjMG0hxoPi96hYlBMukCbyuaQrK+0U410zsXMvllGqKBstqMoCixgiRQaN
KnlAyxvipQYXc3bn1YuM+JRTyw9gWJJdLMWBSicX1qOboMCvpU9nvui0PP0hPsSGzv3dRFv+A4vN
tE4jC1Tjxv/vau5YGtsq0fzkGoMJ1kcLmajFzDplmklRSnj7MtRcy18l3nNuZHmdMVnKBLGhOJs4
hhAWQcuOlD6iWYdP/VRze39GmTlwxcNKFdaTul8wBC8scAtgmfyb2XgVIhDluVgjuNNdoPnUVqis
wv95zglAm8hbwycaTHExG9k7NEYPkIwvARc/2C5CqyV0TrY2i/JtXzMfsglk9m8HbjTWp46YWUZY
djXs3uTIqdnU+M6iKX2syBoDxsO056YnSCIIrzuYIm+OwCzGV1fVcsSy37+Mo44zQMKY5AFmnOzr
swEC4dAGJqZOBt57o24qeACxadHS3OyUmRfrbp+Deghd1Onnhc10Nv+3cVYOLbg9nsnuW0fy1HRb
wlRlZXpmZqm7VFw8VTUbl2POGDgBkYCN38lPIhpNVZUhAFIo4MnApKrpeYfbLgHnxtHJ7B+9ibOR
r4X4bQb6I2G9MAmzIFrToencDoVzkYiy7jox2c+AnjmVgfs+U43NBNeZP7tSuddRIF+WAHN925ms
qhSgYXx/zHCLPORkXZOOy7EJP0InqfNiQ0ylJDJUgNKPNL0CFrmce78xx8Gdmj1pA5SPHpIzNt/s
TXkyeS6OCCayxLm/zuy7AVHmEFoVBs/H7BRJ04BgyleEBl2U9E02RfhARGzaeSWLQLZCSrC8mQQI
qfLzlJFN4b1X1Rqw29UhFkusxyw8sO7qY4hEt8LTgWddxdTu/VD/LxGw9OZmV6gEOsGQD9MUKA1H
k9atEIW72zqDX5juKADegYWkfmTFdgE8WnmVsc2zwK/2OEXqLspeeCd4fokcFPa/QBqasewJ9qGb
EDTYtdqU9RihT0hzgR5VkvcAXINzbhe0Gt/aK0FfPDts9pLuv60eY5gX8QplWgMTFfOJOewPvEWg
pLb+u995XhoKT5KSjPhp88pPH1hypFrCgycN7GUlVPKBkCgbfOD3gSY6tPuYNnw5q1sObAnp0Lky
ZCCIqDxDrfCOqJPjI6BdgZYtTpUjnBYz4fllRvDn0W/M4L6YKcKAuEbBkM433Z1EzjdVUE5VNFTp
0iUMLpQQnumgeG4gyTMT9Io2x26jksR6GcISaQILSuIBVlH9xkvXuBqGBQYCQ6kFiPNGz5URvwZs
xn5RbFLA84JkD3GoE0MIKwKYldYP17DTHqRfo/mBVrrnGeMAvs67qzyJYKuQ67R06wc7imZ+PIur
TePdyZ6F3raOPwUbf+IuGnBCwE39Do5ELwjU126Dr4BnfEF1sZLCCGjGHe2hxeZeCVX+I0rbjpaN
Crv4QlJ3ulKsMHCSJbTP/Kl8U7zm889NyZcRa+HGAsA6ECsDvnGhr3hm13lymWPmE9WZgTeGirUP
H4gQPXwiy7UH/th2l3J7bjTgYggYFEbrzS9ir5OdphLH7o9TISrOyeLPr3AkEtAWbwG8OAkUxX3N
NWi4klWJ6bwCQ8u6pOYVtxurEqyKCU7p3Tf7w/nGR1E75rQ1Ajf/DIMO3I+ECmSTr23VWPfUdWJ8
f4FFN1/8xmNarqHAT1bZA6ROGAWwgBdZSXnYYf8uVd56UAcS5rJLBhugIFeN7VHpVjitzyw6ZEVT
AYFIVoMi2eNa5HbA01kjKI8I1P+aP/xmmI9RAtxkA/twuIFWyW4YCKZK7lNpFUu3p9Eo/X1n/dp0
OHREvloFLb9/goyowzwtUduq1aks/fjB4upqKw2+bxraFv07ZJBa7pSQ12eBcne+hnqcZd8/Vdah
acNy6XmmMF6v5IvY/zKI/2pSDVjHr94mBdkI/AWTRcaxDBQAjUhJM+9eDV1qtkEhq0qxoKx/TFoN
Vgz4FDbY7flWKoF7VuPRmH1v4VhIgDN2rHqayCpb0nqxz5gRjetQ4CPPJI1FvUUc26ULogdSTGOP
OcHJzb6quhhGyWigIDqyjS/vbdGeJ42g3Exu8tOig9Ln/pV7FOrKCqVzyJCzGfWrTPJhAfZPj+2Z
QYpGhCGxLCC8L2tMlM1z3NBddJmnufxCiVzQDFrRtrUiRuSwASmoQrRftfpOL7E3jusDYKcjsxEE
OMwtJ/f8pTHZGiRX+0ritXMPPK8HDrgezFvIcZaIQo89nBDnXEEIwnmYX6mjTe638knz7/L9n6tt
NezYxtDVcODH3fpjxdzO+q769obC6Hu2Q0JoCyeCiMpLZF3O/SArxtFS+spuVO0FWxOZZe3IuMpI
q0e2ZWsVGssFwD+gMzjuU1jjhFA2UYwAWCnl+1/hABEKzNrPVLD9OyPsb8mQDo0IrDfGGeUoEZOH
STq2hDCPRflUCwGDjOSv7KGMKM+x6ziNRH/R6Ifi++WQ3bQJ4XNLVAJqGiYjI9jozSqVE/hPRI+1
vqLB2z67L0/YkPQ2eFEsgcasY/7hmXzuwQfAduHgMdd92bh7nRx1g/dRSekmY02ptJXVfplJq0Bq
mZ2RNY/riApSWo2IA41/qD35Bzokes8liwqBdCfv4lWTm863QTogEtV2UMNE5xLDKiRHROqFVzpX
K7mIjVhwa6cfbMX76O1XeXPJ0esj/GxrMVrIwsDJxPiCogF5w225TaPpcoPGo9l/QI9FFnLzR0BC
Jm2sNOAHJSImQJhOUod+3wKGOOT2NDyRUucOfm11KlX6p1MtU+BSjgvc4q1iRg0CGA8GtXR30auW
2S0SJ50Z9WAfZyqotTSAKg/mpPBLCrYprNW1gbOj1yfh44AVgvwBTmvaP/h9JEvrgPHif0G/GvaN
i5AjrFRs/6JIOHr0bSMGc5HnHZyRVavp29oX462tnx+VUusSXyO/qDoWIo+HGL5heInsGnKhk8qe
nuvkLfMjFPB85xSkM8ZaxRsFKstOCOw/xTew8ApCUJe8SBXPIkAs1IQ4TFP5SYK6uvfgUQip82Bk
Gog92+67RticPNPDmQ9KCR+akoE+fsnk6zHiwmN7pfPGj1h1m8Uk377bO+xAk8I61j862XlCZwnq
Tgc5TI0bro4s5SXsSlggGd1LzWanGpywsvTnT5yRlRmyiN2QdaC5n2MO9eNQ3xgekEa6iBU7hvBY
QKDvudL5IQXIlOCZgKQtuYepOs5C8PDO0Yr3ETpFBn8dgvo+dzK5qSjESvSEFcrNwYGwmzgtadEX
idX10Oipe55lOLG4Qx28c4BZc6VQIj/KH4gZueF7GTOC9E1icC2Pmr5+Ca6V7Wc/q9LmfvBp7l2F
8X82Y8iAkqvLaZlPy3svo+DVkTJ3o7Tnm+UzIQAtfAmuxrc1US9TSLrRFIofMRKbDykXCPko7+S5
LMfXHCSuuRTxsSU5rRj9eCiOjYeAxHQj2Xyz/qM96zsYCU21p0YX6VPf9NrlY0PMleMt/PNcAyWw
JtjUNUVCU/fxq+mT/HaiN5S8BnVnGeWTkoKtW6AJNJXieDnTb+Tm06JNWmIYkDlEIlV30YvafEWf
AeyXe6umI0sJ5XfJDx1RZGM8prqRDuG1vkb3/FY+Sm+n57LapD8rtlIIDqLjT2q/ZR7fzgzLBO18
d6f0w9x6y8NArwP6j9qHR+hkrVOOXFnSjarj8tcIUNLXiA6IaKc9tsqMIeUkA+ZTFG5C4iwS8rvu
djTIYbwmvpfju7fzQMspBxTRYW2N6WoRUicOQDnR9XncUPUnBcv9fe20V0uMOT65udoOYqcf6XEe
X/eQt02X4j9KiKqnbr/jofpDPVp+X8SboTInijdRiQz+0dnvNLkhXPGbFjmOLrv/xfq/Qh12E9cZ
oPw36Yxr6NaP0Bw946ZrvnIEjrlFULH2M4WtTvDV5aXr/wn8hcM4t2W+THo0UX2xGf+iSvdowjZ1
VXKP+cZEZwGv/7gjmkjqTIelIjedRDtmr5CUE6U+A96zTq6n6z/WtHcQWmzFpddLL5zuvyDVvU5R
smQQm1V5QcpUegeDoyQdy8l8nqMINNZGTcJztS0ipFwkkAxFO/+IG6JIiLMYW8HA7WiHl2Cverld
Z7Vr+9x9IHFtXUIlYbD7V8i9TsCEneo1KinxQU3IeWjTjeFidIun52d6Yg2QpbF+9Kffmm614Ihx
Mum8xlEEGNrX7N0dvLKPsYQluoCApYPphheonOwzHw+nYIFBmIiIzkbKgCvg5evJlnmndM78QFkm
l9z9vbFSU4FuEc8WjlBmJ9z1tJB6UTCEQS0huL1uYg3wAoQqbC7oAjpAP/4x5Si2jvAX1muTntzh
528O+ZxUlEptC4oy0e1YwBmta6lRryxgyR8ce/ewLgt3Z0MCI9Hx0s3EnUbVdO3DuqQi4CebB/5D
mJPA0Kj99wYRj99+xfw2S0u+28suSOMjBy2opwXqTHJbZOs9cCgbrWzlHAQy99UPKB6E2H59EQd2
Qbbp0fmMzv9zxBfIavOi3LX+gIYuRbfcnBlADAaALgcjYMdqs/MF9CNNTGb5ig+PaqK9T4aFodHd
G2xoj3jkpwFdffSN5EPkt8h0Rl79i6ar/RZhzW/N2HsqlT09kkjNWYLokry6JerX1iAb2x6RcSYZ
H9BXC1ufTnJh6PPsTEXCHTI+QAcc5a+i0hcKVG3/mdK1uLLTxbOCJTBgjiHsEZKV+shgC3sYLsYa
pVLtkB/h/2TmhsijwzG/BpabaKYdp0v+jO52Qgy0iqqo5yAcsD2kAhcYJOii3UoMwGhHXpGwTLd0
QnqJgidsvCveONANZmV3bfTYR3RSYEpQmO0VcPhLNHxqbOK6BY5xjylgu03xLbSQwE5EgSeuql/9
21I4apscV1KfPdkaCuYY8SiE4geRCvlxZbSiy87tPL90neELDv1xL7jXlkltyUOwtCpKh0Z0shJ/
5MYwVCAG3RMrKUZH6Omya7zS8MavjmAPGV06uM+Msa/EGabvZVpLV66jJUsm4s1Pc5ryTR1/0GUl
XpNGHM0BDwEz/NYoxL0lx7UcEBtfmZfM+Ck0lQVFnaOMthvH4NOYZQkHA43Tl4uexDHh+HUzBLZv
uAJaGUF/R/LtD0+9N7xmazuGByDigb+9Ol6yuumiv5aQkPz/8qmUqCYyxGIhNCANqp7nJUFCwxsL
fN3XEEdgbzTo0nOFbOGKSGK7bgtb3mLAIThnlQ2qbNz0bBRNO8aKrqwBaF8tEXMj5SH9sVMYcuxe
9ah2VspATl/qHL7aQDvtFdxKEG5VM+zINzZn78oRYDj9RiblHBNyqhfq3LaVPa5CaLmR+cfvYdrW
Mcx/w2d/vnODgoT2idbczTbOLrZ9n+tvqe5zRi0N4MaTR03k0Dz++XL+xiJb0MsiWE85vm0aYZgb
d5HbTdMnv5ComAZvdg720gi+3PRyAZXz1FT0meRxxltIkUGzlMdAUHtXzTtzTifhw/xfSHd9Mkoq
iNrRQdBvn/n870eWlIapXCuVtpDMrd1fNEusYdDjx8aXg6djSRaPuHDG4nZGfJa3f4eTpgxMaWRU
Vjcdq9vmAhSs2dvJgZFPapmvqfTA/3huui9g3V3o9WIPzsk3anyU+XPVJ/mmqTPXprSCdrMjkQ3a
CwBQYqX6cMuKKQ4vi0CciGD+nzz34COOCycRjHvOBf2j5ytRnaU0/b7HvWGSTqHNHNLUB8RabGVr
vdFIrNqe5jI7Ptg9xbPDDBhOvaqSVeMmpQmaYhZige8YqvossN07WPI+44eDneNG0Wf0wyQ779cV
OSX0SDOw9LKvKLRRN0QlXfyLv449S0Mdhy+ZwjjvbD69uLU8wyCZ1UVGCry9OCkSf8WAc6Ok37xT
JbJnc50dZITaoFsF30vFE1rxiJcUqasycR3z1Ng2mXIxBzH88nFuSlaUZ5FMP8kymatEDKYA0gwm
i8XueRaee/jhGgjSBh3ZM+mf3E/83WsAk0Upw3d/tncCb5isLzgSk4gs/6vZ5rTinJWhTDERt+hA
G068++Tlu2o1QK8ujLAucGOdprbNHN8VeAekq8LTG98dY0cjk/Kbh8te7fm/NBZmruuIAeg6Mr3g
V3gR6xbAAfrA7rTAwqPY4XTEolTQ5eOJ47ncHyiK3bbW0HEh3dbvq8qkBun5jbIO7KUfqH7qnWT5
x9NB4xKv7bMc6oqjOXPtV//B625lqVcO7HfetnPOL6xuj53+FKUda/CDrOLWhDj9AeBoGn2mJELk
cEA+nHGEzNtcske4i62uII+Y52GYu3nORKv5A+W3fBZzpsaY/e8Gl3ZmGZGlbegpKaEe6p8fxNFy
S0eMArwWRkj8y7W2dmTPW2IyVdKVVDqBitAhqjuQKZi61ON1T8rpGLXNBFK0lCXVDMtGkmT0+Gdg
2wK9GopKQugvdIlnEialoV7LbbYSCwwiQkc0wQpnn24z4zvYOo9BAeHXg2lBkfb1qb84Doi0iQ/8
yWcRfnRWspCvVKBQfq0fMiZM8OtBkrpsAwq4+h5Jw1d3HoDfCPYozB7xZGQvpIUsKbGRo5Eiivit
qv4Kd4MqmC11mofJaKC7JoPg+mM/PmTPBrQmgMmGBAlTbTspZScuU6t9bgi0kYtiItvRY8Xm0H6H
KG8vvVqFQJP/yEof4BhAM6upjCTIQNDAHBXI0KeVnrwiGJaSxaPDlXJ7iD82EGwReWofn4AxnXSp
5NCXxFpJtBtNoh7XkApxUrLZAH92vXwBdjlrQsMjlyKaktT9e+KJgwspr5mF+bcpm7/ekacPU0R5
3nPyC79h6XSWxhAnhMa94178bT0WQb+zMGCnjp5fU+eSqWQY/qjpX/XqTORxoFZZw6PO+1iG3Dpg
m5cPoxYLeg7OAihm2p6QJzqtFMBLHiyc/Elk5K3F1zNf8lxwHLkIUMS1E2UQF4MP4qmhby+0IKIT
zzam/9ES1elmX6skgw70U/7EH9Hlfb41WKKbmiOE4snwRNRNa0M82KjbfJ2slhPnVUu4qLhCRD4W
Vw9P8Z0u0lPfe40r0tkyRxaZiyhS4IeRUempJx0gGkBw/MFYrRLJlzIjP6MpSrsLpsZsI/cSGhP2
S2SLM+EDuXpPrxaEHIfpVOdQrGf0mKnwMM7jtKygs526r+A0Gzfl4eA31azJhEowUSrm2JJhw9ff
QXu/h2cHKpX0EHCFjkA13ltEScs3izjrufe3FqlVOPqnERVY9LMfpXzEtd5c5BjxKul5dmWxkwAl
DKKeY3m50E0TYSV5tCO1qRKjRfS3W+pSwZo0Yu2UIohxMHlSu6tKQBPVwfUqZr9J2xmDQ17ow1J0
ZvFxEZ3M4sc9ZssScck+oym8pjAOtBDa8wPUc4DnIr69hCUV5R2rcIdmcuOeubcxUWHodl2VvWop
n3JviewpVo6a4pqMToCgPvTNPxTapDyJagwUEn26ubIrIORQrb3tkG6NdiYFnlJ5Sf74toQoZi52
BsEv51odEp6PViu2wVPW63f1CkuK1K4wJml2cUX9+EdErSPDFerfwTHFIIWA/aCca93C9mg9NQEs
4SEiFuP72z11zwD4G7ZC/VFBQwHvNbpe2JqjzORIFOlVr9TNTzibTydxqqEZJ75R7QAoMK3S4fgc
wn5LcFZc/dHlIokOdWOvm2MU/t5m0SIkPYnm0vjgtOVt0tq+W3u3j/zFFVzOBRhExbhr50AhgKrr
oCgWoxkOO888ja1vH+TEvk93UDJw4Dy+YspuL6w3eHFHvHzyv5bvCX4OFYhVyciabQc/5CUH33F9
9QsZ/OHbhykz/40kYJRmhjc3cnhsv7xQTStyIjxbnpk3i1SjDNhUEx3msgTSdSOMl1W67hVIa6FZ
79c7bfmhOuKldVw7NzniE0aeQBupcq0254wXrRIMp3V2P2d26FZn+NLXyvkSv9QtpDAtpHJ3qmFC
BJIbZtM05yAVfmsQYVXnOBc8yiZ+9aHqFy7WTtLVx99Yniof6+bUx+SI7SF86mHKnxgmHD6NxlYu
ZGZZblPs4AIXazBvUCarp/OCQZSDyHhF0hMXugRRDWMfOoG0S4J/9d/InhDN8iEZhsW+n06pL5lo
tKIKbfXMO5C6NIDOik4p6QAhUqCRUayeaPUGsbZIQzF7i8aVQ1cuYQTzgzTtYaELYqyrsqM2Q/6X
IPWb9pKCLXXHrTxLJ3lX5k9ltJMCoS1LaiUrKtsO6LyP83Coi9uJ/y3Tut4DamHs222Dsh6OV940
2WbVxZyD8/gZ03rTZMVAWKjrXmQ1EW5W7G5AX4sBDq6P8Q1F7+Su/sq0iwhC6wz38IzHCzSiSD9k
75iWIJ8asAymsUt5aSBODkISZUNa64IFo1W8XcToPmDeGc+36nGAAK4kNW/62vVWPwhs8WHYmedR
EnTpcls9r9x+EavdwyfWfMrvZbf8f7qxo/R/fLzRSbg7+pMJdHOBUo1FgaNPthL7O8Eh1EjR0VAf
tjhGkGa6PnO3YicW/OL8H5fr2/Rd00p9upHt3Fhn0GG7IxH8lpP/hk+px03YTwHMfSU4w/FsrcP9
gTLPbkCpHN7WbeXTP5JacWVeFfxz8FMCcE7RG9hw/0mPTaYSz+DKkGlUcYGdCqKy82lXNVwMdiYu
BpXTFsBDxPji8ivqs8NrV6APlKZLFJ8hQqtT3nOE/0ZH7gwWYpFsCIib7NrOCPHmOOgeVSlPY0b6
y2Q6rFkMhMxzHVymKI6lGmVZpGRRmfjSaPUATSA2u804bBY1UGN4pwPfMxF+tv/9FVSkYpkr/rGf
N65aMvun8Pb6GK8i5UMt7mCFDBIfcg8gFTl5gdzr9vitKe2kYPuEr+x3DZzExd5sX/tyzPQUeDLQ
HVfKt6/3Pf4OeAxd0A5C8tJHJ52V6bBqxoUtIQBs50A0Ou+jvHqSt//6gJxWq5EZLEtnHHDZ+cZh
ooSQgf5uq+0zX8c9W87oQkbM2BKCk7HcR4QTfdSEYBrz6QHtzmdK3Vr15dvQaUA2Jx7jCSvwCvBy
EmnJL++RCWcchQWhIi4Dfw4BdJNxF1cvOJpTl6GNvQ3SqumPhHwmnUBGTFRPX+aeIiUbvmyczI42
bJyW1SaRbliLX6tV2xn+xfw5H3wBSvNoLDGOX3G41CuTRNoFGC1+tgEA8KqCjR5HQJmdPZd3CjD1
fm4rnSAOhx7fuZJc/zOILpbv2hgevwy8affPCabX0qJdmwH4KqISUWp52tqzqbNISjZKFU2E9rqg
QZPpcJUMzpBJJSGsHvwg4NQ+eoz6BkjOqR4jMP5hFBZyJxMzftyL6U+5vtjNQQKv1tT2qvkSJshz
bWicB/AApS3B8/f86UnFF12F/0mtst+RE6fjjCNFj/pC20eOakb3WJX0ql8WWGQEnzhCXfpBQoOS
oUyzhwGUdVrinURk6LjoOJmt9e9ac1+GP0drRPM0X/hoCwqAF+ny6K3qIAIccIx57udK30sKzJ0L
Kd4BzwoR5XPskiN9SfQzFT64HoOgTzTCvmYk8xXkN2Be7Jzcld9Yttv9FnA1XuVhl323HjlTexlt
2WRUiFKp5hgjy+UfFP2Sow5WS3zQR6M6vXrFK2je2PooXL1ujQhbV1PbVsWD6gvqTPbM0q5lv7F/
flH16WQCyaWQMI0rrETAaO8Mhsm7wyZERLo1UjFYo1GD7jG5CwDj4Z7X3LiSKYAKJ756o1c4T3va
R9YCzlWvaEldF1GeGbs+u0Pat52BSkgVEphulydrjUmRLbjLo6oUapy729brijWcZa3nrIO9ZJuJ
bmINRM6mc94vxpzC9KPRWjFnZVyFM/6WFjpJMlkz8IqC1dwn+rTr1hO5azXo9T0LU8WREftrK7uZ
euibxcLAgxlo+ITgQY/yenvPdMUDSSio/kGZi1t0JLPjfU38YYe6ao3ZDSfrUp5w2xh27Km8RoZA
dlSmdeqnqmORTmtOEi0QKI/sboFeI1XwOBZBpnEZrWPdJDcRBJQ6UclC7ARrFobzT5D5W1qQvSea
NDiNWyUtu7eYitAXA4mV/zSBM9p7n/Gs9wz9ufCBhsv0gTd48zP0u5s4Lxwpds6O547YTXhIAKKT
df+BiZZsXwxcq7aZbvfIwgHYSYDM4RHz4/89VXdTjrh5XlddHmFUD5jGhCWUMasUoUpQZ9T/41mY
8YHbDdTnTBTPQMgLAdXDUqmW0hKNqyeeNtR/Fhm/rw5kMCQt7sd3y5dEZOmAw0+lx3lMiGn3erG+
UcYOtUjZPXPpD7McXX2fLSzE+wjFdS8aE3c8j9HUincLIIre1Or/k7KYNo7g72om0uP+1j18CnVi
ktjqk+kirDAq6udA/r001ro8Lortq4xucxhyK30/JMrA3zlB7+p27uInOjk6Kf5jLA/wSZ9014vs
a1xDBaFxteQ4Qa2WuOLzYMzR0+NiUA6Q/7oVoeUfeUj46yQavANq7wmS7oeKle5asR5z7Sn2qbIW
YZ9Fn/SKx9gMPVejERzlyJOnQEQkkmRQmMR1dvdz7lLabNsZNgjkHjSCRM1aKT+QBUTr+6yqc2nP
TNEpdk0PGblefduJJCDCrFPQdpNX7egpCrvjOAo7UaOf5CIL8zoTJeHu86chjL2PTg3P9u4wIeCd
DHwwpWn24IX8l2wsb/IgZ9Uvh1HaMic7knpuwMaeZTgxohvhfA1NVrOsQIU7/kX4WU0S+tmZWHd2
NJOM9RLVCUUZjOMHK5w91rQ2xhd8D7jwCkMyTXRR3QMqdkdqlTnQJeILS7cD47noHkLzVEbAT9Rv
0gcJxRI2NFBmcpk43hAz3G74/ptAIE9n4/W9Yz1/pMTZlC+MGQFBbVO295kLTxv4qULDlXUa/dBg
NrQJF/L2H1DEImGTqDcO9iAWl1vakQ0yu+A8AqFNJE9NV5bMrbij/bGmmxZb4pRdzDLTe4cIvbel
Y/Hdx1HUU6obuCdSTOkaBKL8LfNaCrneaTlCTLGGuM+D5edWv42MMe40e6Kq0tdwsNGSjURkywO5
VlFZyAsKnR/Cn3jFvjDqE+ZlTbL/BDJ6bSWIfh0MlGnjaMAs2PuKvN+lovupQFS/BrdRto3W3hK8
gb4fSaAs1owXd+rOE3QhCCE0lfNA7WpNQr6g5hBeSUakTdRIwledi+/iaz025St+qWHllxWricT8
u4tzMANRgO0yMndWqTF5UIX5vMfSJE98+JrQNJEgPwLjA4JfCBPzOZ0UfUl0xjJmhpgw9uwDCya1
MhVB2JNTiGptrPd84HO6uytNIv1NBAr/FivukRpCuMWUvAzcva08P8A9TlH26WKbJFhDxygDqMx/
5jY8vl9yerFF7EzjrPuzIr4SGzSKPYMKaKdrLQS1qGVzLtTotXvfuQtnsP49/mR2UCH5mxvcOmOU
wktOagI1qOC6xmtJiACQnQ9K0boVFFC1ULB1hKSG4zqRkNoBtu5IzzY++64sj0RCSyaGdGcqVnkD
XumJ1UdZRPpqDABnVTYlP9s2Kpuvw9t69DIHKWPNhuDJzyZhETMsLLDsreoG7Jrr9IvdVov+VIj4
diLLlM7tOPQfZMpq7sVM0U/hyEwulF1GKXERMbv6lV/9V7ocqFVIOAQ4yuPfufHrXhlNvwCErvwT
8owDYAi0VjreeSvg12Mw/Pc/dLkhvb96iI7hbDcPJLWl7BKH4nsnrN8mNVBRfkHtEQDXHN7DXkr+
EZkkhP3JWfLtne6IaY8lZY0V349mO09ubbL193/ZgYZjVsJsRBqgA+vb+Brn35nZ5DZJJtBoP7TY
KOGsLFa14arlkjv1ZgXyFqe98MYAbO5oTFAqmLaYIHBj6S0m78MSgfHW4jUC45ZnkzZ92041n7zv
/P/17sYgcnY6PcCuGCkiowMEGWlhvgm7165975nqgN8z7VI3KQVARmP3ofQrHO0vXaYJqc58Ovez
hwFKCHM1+opqmoucJ8PFTn+NoPbbnixVHp9JDJ9Mu+bKQVPOL2EAGCd60BtqHRBsA2yIKx046NeC
JjoJPhDD+7MFvJ9S3UFXB7iAcjoXQ5xJMUogFPK3T8QJ7j8l53uEqD1jrKjucBSVyHFZl0zZlGuA
sd2L+aVIvgLWCMwqPN5WyRWsno2lWteyoYSE+gBWB5yNBzJ8T928xDy9Jc6td0qbvauar7soZ4FY
Kbb4QpvSA2Ey/NTQP7vT/FxmazVtFIaf32wb6fDeSnMzfSuT/MaZl7UcWT+LXSWdkeZ8xldYPQrc
pjYqEDF7kfNqwL8sEOcLj4Oa8OgdqHAVaPUUte1ozxZTFSHpmztIKxoebibsDRhdPOen29ConaBG
Ut8wQZT+yf05O/bxJxq+FXqigI9jdZMYaB0hIEzTgtgrENHrORvTZMeu5naJgG0jIdEj+JN7RBdc
+hs3yjHPVHXyvtGQ6khPP1Jh+tiTt/RzGu1Qv2POeMTDjHh+6dffGvr+5VZWk3rrat0W1K91wAKp
F+xgUkTn7rlLyyk/ykr7Dzr6/kkdQKrYc7VpyXn2KaUCuQtDMSq2UcvwB29hZz9v8voNT0VfHqMg
MeqXC8bWPSzh80Bw3LdzFZdKZHC1dfiSLLKXL+XvWIRo6BkGifNuZhvCGL5+nNRw+l9awMgXpI8P
WAWFxEx1zZriTmqF6S4JJUyJyzHrA4Vipx4O6XeuPJp6aHw4Pqsz0+08Qg+pFnLsTdkcWc0PTmnp
wheLh5HKJX7xPYsEauc/m4Q9Y81SH/Rn/pyuOXO60UF584YxRQT0Ut28dlYOzq3qKtpPEFiMs60u
aKnuNPMZLtyRuhLOkvMLdijAjBbHpNEhXx2GZFAurWQKMX00bFt5rVwqs/w1OgFBTilrqYwFFvcM
7JVf+odUO8NSCgaokjdZMbvqCwBZfxtNyTO928UtX+pQNpigAhVmElFzejvjL4mEi2ZCrBD5qx2B
gw4R2sUzxmMCOfuG8HIH/KUYAZjN4ABuxra5SIgWG6kIoDP3VcaVU2LEbVwdePWHG5x6/EvmrZiy
128ecY6U8vxa/S599hqoNl5Oqn/q34yp38338lOClQ3vNyuEVRyJwuQTv1TgSP39/9Ni1gBiXL5G
lNOJwcwB0ExdwhdcurZptaTQJbLN358qB5lYbGwgogmwoN/8U34TU7NSFum1rER+nEx1TfXJoz45
aQOBlkNichRSO1LuWVQheVWRyQL7MugoyFeY5kBzwT+faogQOBA6CxfwiS4+xWeDYYa0Zkub9T30
JXHx4yYqKIi3KdyvSZGGc7/FXM7kozId+dVbSobZsSsAAHOYJP6W3TYVIIQ1Iq+zyYW7eQ8yj1hH
arRV5m86lXX2/d9z4afYPta87sEX7Enm4yWdjgo8zQaItVaZGvOZrcFiZkw7CIMOxiEmC78NJj5Z
xJFVEIHg1JouTqI8LaKk5Ert7nTA3EWthjx/ATbfGZg/IK6783czdlYbuT42HLaFO4ZxxRPM4+i0
oay30w6IZqcUoqqvqcYguaK/vxv3mFtdQKvN5Z+S2n8hMlehQOhjDjVdASsbX3t/Z0zQjePRCiRE
nvwQqEyD/BGNc6HE4EjHCMY75qzkOaWiPu6IQNDrKFmnDZoU1i/ggjyoanAURFFskdaP3T7B0z+U
cn2dBrGvp7XSV/kFYZ0oEwEbyZsXPL+T7zwNXdhWQ5kGZgvV3NuInMkVKL84sqVWBIJyn5IjZB7o
cv1/mbpw7nXSIM2udZEzRJonhUd5Lk2wmhZm20Qd/bPd/RGeQOS8UV3HAqvcnpK/IsUWTY+LowR9
Fvwy/06Tiv4LjmK/kKO+1+LhkpoF40eDsuDMEy5SVxgnE0HRxI0kNIMKPZWAS2ysv1o1HVBtx1tD
pYPyrtadrcZt40GSw9t6ZJ8//FIT3Yypo+aGodE7ItrDouXkWhvZyRvp3wVXHeyVdm8weD39mpop
pvSJ1CzbZ/QKcoWfP+BWyAHuglWuy3eXRBQKGjc/Kf4OCAKy9ZdWb3ltGeOMp6X+c+urrMfiimnj
kvcoe2FonWl+BFPCDpDzpzexAErI1xecqv7ob7acYnmvBRKjb29dGmxd3P2j2M4Ezx5itxUzjwly
6ABOF91h6e86bkVJvfg2OsH8Xgqr4SU3iLQqyOwTy+yVnOKhGrcr2o5Dm7P8vH8GKr4NbulKDZ3d
2rhzNfFs57C2cnBjX8HGH5Xi55VTYBn38tFBbigFJz2FQQoVW9EeGpZ1J+sYrc+kdXMJ7uYg+RSN
FdBPVzbk/BU/aKeHpOTAXYZ5+HC4cTtWgJq0+mSJ8U2sqovwIq9dOayeQijjNGsFEykb/f+AqdAy
bDRBMlRjJ9uDp6VCYlAsC+HP1WhUC4vnxufn3v+g+qxxvY4n0oTPOx737vmiYv+3rxs9bg3HmFEw
PSHgOThD7GH//FoNi5NjVD0nHEYv3lf7peHfdgapxzur2XCTVLZIIFfNWS74P4jCLTIIq4t6oER3
Up9bDdXbKJQPD+KgYU2Kvv8yMvG637SQ8JWXlTAOnnRWZsnEtyPYOotEQC9izceE05vt/9FyzZ9a
anBfg40DR6BGSmUQmXsNjcas1vL7ju050xX12Lc/ks2GyROEkOqdU9Cl6+sWt6r0sqVyJM8cvzjs
z7bF7swlv2ZU8/8RaFCvbROLWgVvzXCI44WBp6rPsuzWMmD09L5Bbf34a897PQ292EKF/rCsHkSh
GEd3/5TDh09XdJsC7HGsILR8d5wtKFIMWkR+tA+J5V6iJ9s/Tu4bgDJWgfmdlSn/pK6YPKX32jsC
4G+WZ76PV082MEMzoEVDVOmaI8/o+bajES3Cf8FvRWmIC7J6I2tzxDyHE3Re1+IE1eVJiEAHxixD
xe2NL1O+Qoz7T/09sFD9D3BY+w2e9arABxnQgVwe0tjfOVsd28Xp1VFaGNbACZEL8SEums2YnkLM
HPgyNYDBzYe0BTEBZolJhGg8i4Y63PlfTyCFzFIg1D19EHjqly/8chAKylc398j6ctCa0euPmLFB
cKBsil4Zv0kYlVZsqCAvhLr/oPUIJUeDvFGBqCKW1X73xNuDv3IFYRyNr22nBsURG6g8hhv81S6A
YNRj8a1T9vq8QID7nR8uIIpx+GC+Ej36Ddh0/zSUihgmFFejeOpUfKnLbhdy9NlW+dOTajAhRMcU
8ztvy5Gp6zvjrkMPFCT/gDN9YMqLDVPAr+4ZbAmGNZT/NE1Sw8X/pzzdTsxAVgKOskQ95x/orl4W
vAfpz2XWdxlkBI929N1grgxbLVmSFnjqgwybqlDDDpWNOWvUx4yh0IYm9yUVR/YxN48bx3nkH9ZZ
OYJlpKskqb58sv2aJ9UPySnW6RuWJYlmEU8YxwW7uGoEHOZsUWCbcn1ptWmyRDAmgwbNQm2j2rkm
YynnMs+/h2yHSpRkpE/hn3UhUSwvOZVVt8oAZ3ODAH5KjTgBU5Dfru5ERHkxSOXMWe/XkJivU9wI
pW6C9bOy9xMEVmoofBLfGXHEw/qQm2ITn/BgEI4GeyZly8b20WGO0sLggL1BSOyGKiuTESb/rjbX
/l04C7NO7Z3lV6YnhBUZkb7qAZ7b2PpYLbbJ9hrrufPqdM3avGImcthz62Og2/XXJCLiKm17HVg6
+Wde7KkkeMKDmiAn2nXhS/K1KF4zqkFSViFknhbq4Sydhn9IdlJSnV9Sy6riMDArxn9KCtO3hQn7
/hQ5dDwQG9SpfIdosOQpLqqVfbgsnXYK/fQSb0sb6hfSvYQWlS3/nV+elWMc5hXsI8ODnO5Zhu6W
TOKnEZmgXGSen8+NBcZCsayGC2TPVDYVwQPnj1qJIjOQGecqvXPipsKmFDrOswzvfIqt1avu19Hl
kuZmpM77pR3vPIu5AigzR/wyZs6ceVbH9gddLAO9HumCzENH4VAWahETaKPtYI7vl/+LpvBDBZqA
H51fRAa0X+FNu8HxV9IgiHgRRMx4778U5S07Bxzpzxw2zjbx/bfrWvipfAts0nnNmcXp4c7cB4cd
H74CuGk2xAfhn5+cjWENmX4ADzuDv/748MIM1zDHBmiXnIgq66aWJydFLgST//0Oo8VuQQPmuHdm
znIgRwfVet4iIgka41oMWnWQazEAkQhnCDNabbWZ9ZIYdwMf7697a/sMe7sXwo+wJhZym6pwo5GA
T+pcQcV/3j1mkM68QGyOnthgrx6FVqqRHsoEpDpYgRjkeZJ2+DE55qG7TVihNnd5h5sgIU1fIgdl
X46g78cranyxqNibionmX1S3tH03d0ULbVJMUQhSL7rDmy9tmjbwYgGKVNuPakIEgLlT7kXrqZ0y
4/FVjAufS9toTjBLJU/eijGq3QNWAEF8k5acGIuElI45SiSdzQKcNhZ3hSGHvBbZ+dvT+e9X+xHl
E9D8z3I1HgJgWim4pS7+jYy2kPoOsP+w0ONd7/DQhZKglSNrRisPVKASqxxfyKtIkJWAD5feSsxQ
hQQkSghmUZheprAqRRCt7mBicgRcit7NZQTdSBOW0S/wv/A2TZ+d2rr3NknfV7h+2XmgdAASubMb
xLYP5vEG1VlZqStt4r2M8vCO6R5whFobXTjfteqy5IyKMKLXGD2Z/MMAMCDL5E/DY37bWfQCePCY
UqAIOq8aptd2RjCOW9MfluIcI0ZL0JuBwJKemjHkuje4sBPrN7OjGmyzdeWjCDT30DGapZHKNieP
lj8gqyAuTSyTAhGexTErAAJsJYcGlGeYBHI+kAxX44Yb5paDjRVkx03JB77mGkK3hX2cLYRAWIar
2Ss7Wb1254SzVe8v42bJo3Og/ZqiW+pGgNoJEHs70OGMCGt1nziPXK3TtL9N5uK9SGPBiHF4jnmM
zCd8ohIXBLQhqiF1snS/wRMmlP0AWMOt123RA3O41MJ0zarXxSwGGlOICIwWzHptWU082O6WYc40
89sp9ZLi2E6Sy1lwC41i3jCgu4BkdI67jR7vbg4sf2TMCT6Ye5LIL8EH7FuzVgFFHCrcROu+lMX5
BKYUjIWD91k4v26g2KcUpkogBTN17J1OrU9b4l9XSRq04igGxWIOhIq06q1kEfzmzIpbDnPwAuEs
PnY7Dwaowm8wdn0eT+3w3C6CA+MR3NMT5hG1ybGLZvTthi2/ZpC/C01XWPFD1ZUJqaG5na2ULl8w
0WaOkRrTfJB5K8vhrSboT/y+Q7w+piaMxmXGFCWd3xyw5tpHrCCMeFG9rEK8XUlOeSQsTDu+PUpe
PGN3oeD+o0sqYPPH7Q2/UeYcVAEGqnk1906XjpdocMcNt+BcAvWB5bqbD9Sf4IJYrOv2fvXP3hUr
PkXnsSPiLFX5j3xw5cHXeBew5AT5nhN1iiq879U7taJYmoaBam3/FuVgXueXwsybe6gN9m7GD5TM
PPw/Soq7uwJ/D8GlU21GzV7hUVNKay4+44SkAPbhGUFXQpHsj/T22OkehIVBAvui7IiF3Hno83HL
f+ov9hAfhkpV5e9Y7eYUySv4dj26wyGbM5ddMaWKt1BP6aFNEjhEnEIK7jIUXrYBVEGN5KfdiGNa
KfR86aZDF99KF3jkHWSKFyQo+t8YbEqY/v/L05WMXPqNBlo/DpsdcgGvdTBIVcGg2XK5xRo6/tNa
i0+KddfnJnuDrVTwanYhUrv/Vp6Kl31N3ufQQJ7qLSXEmU0fuw3HoIuADp83V7l8JpVD3q9gA6P5
ZZNav1IphN48EGHTEVzAsNXT5UtSWDiYXkPw0ybXjfu9ogD01zajlnH+Du6VDwga0bcSYg0MID/M
SKwdOpYwXEfUPJgjWDUmU4aAUftnsxUqvMlIlB91tHeHhcAznS1hPS0QdbWavtNzoWQwgG5PU999
x28s4+FTWNAPoXF1+GhJ7svcKpE31FGNbkRoPb88dz3D10OdUnl5q9y/RNGHRgw7qPY7ZQ4Nqj2n
fAb18UsbXMSScRw026y5n7HUf3eVikwZTJ5gGq3NivFGQc8ewhC1I1Dm2p11J9AVx12cLG0c5Xlz
yhs0fo39/2j681efD2FYsfiCQEYsHbAHuoBlGAKjQtbauyO3csm7P79x4ibA+VYnykS/MDyna8xc
U+qnSHq6PFLzZlFGTA1UyzER+dzcliM2GGQ/qsuJcgwCuCRfiMJycevuKnswpeO9vD6Ro/8sLrvl
13D4HGQ1mxPsfQ8vBSYX0WinjC5aebBcsxomaa2OJCZe1WXi1noX8/WR6AhpiLcMAeCTVrfZH0xp
qYMFrWHP0LI6IrSpqI4IUNhMjhbo8sbBCsbu6IDY8ICo4LcXyDbhj6l9ias/ibnhnFC2faYhdYEJ
1fWdpiPrVflZWazLssVvx6gnB7D5Fp3viwOlqk4uR2GNekUdGCAMQayG9C3GzZIYytjq4qvtlmps
OLqnb2JfGBHyNhM5UrFmiSB3uv+m08DsDgJ1VP80LWdFXdZq0On4iomKwK1vb666gL/jKZMyjPjb
OudLC91cJ9MIcmJH+cUf1ecaO+Tvz/f1jz85naM/dLb6T7Vs76lVfpCHVwSK74L/Gl7p6cCalC8R
5ssoELavNrplSlGb7nLZKp13VJpQwow8GHzQA9LYCf3kG25+DCUz7jPDsyha1d/X5xkKSpaWT5QM
CI+zLlvoLntFEZ2yc6kAcPh85bWm50eXfVXIT/rJtLzI9I1Ii6efgcr9T5RT6WX7fqgiXjmmBtTc
SOgf5WvO6v0xY8bVcCM5n0WTU6mwWNIlcBeU9fhOJTK8VBtn4puvfIFfP8iDtkcPwOfa4WqnKkoZ
8ESW+b9q8jI07h1j960z0Fiv9jDCMP7ks6xeOCr3VMlBwsG8ywcmhmbdc9QcZOcZnlACQ0mi+Jr2
qTqCABG+1rjJ1Xj8gKoOzqTzfnOIBQSMKwwMn/lSfrjiV+yUzrH8W6cPcFhJI2fnLohHMn2mVdDg
r0X9Qq0Ftwv1vcxBnQyq//3rF3xL5t2M0VD/tgSVU3t6+G3aFwpQS62QE8o4FY5UoGIYirtg+DWg
J5tVVbwx5+qKroSgGlDF3XxeUGrHEzxWYUezowTpfCxabclhwRiYp2jJTZWht24gbQWsxmMepm3E
z4N1Kk8CGKWXZgrhX3lC4aePASumbzcNeW0D0noDhPN07MWYZ+/spWIPTM7MftDIEhIRz3molhCn
Xiy76em1odZ276KTuLVqN1UVOoLgAc/DKuFoLkcgoTnPYyHksbeEqL/Xp24cWZBc2RyOkvlDvefK
qjoJfT9Moc511gDWm9Fj+A41aM2XTBQF0eB9cMrsWCfeD3gJGseZtzuWT86mnxMBeN5YR89FFSdg
3rHuhNNPJWgKcHJ8L551yVoYqZNoiLygsUh7kxMbdin8UQxLMCNtxYdoG2t7I6/aHGPds959kaq5
gkaekAnDp22mIFfw8I/AeVd6E+nYczRshl2aI4Oe1tn+XTG3wETCrWbFajUZrbzhS4kyyevQ51MH
NygKewdO3X2mTAoIM6RL/940fT+Ox1IgHl2Towi/UozX3f/mQBznjQYN6ajd6+utB4h9k9Z7QO6y
DCB/vbWBWytCsFfdgKlgm6MLGz6qMFNNvHd99ZZINczO9y5gPrKE+zBYR52t2MFUy6D4mz6nn92N
kgwAn3cijmeESF55EnNEUm6pgSwqVEYmQoL0pyM6BOVPsLDTuY0+5fEbr1bVJ6JQzmNjOMYGPDxh
vqmu9PNhE87iRdqg3vI87o555F29wnKSAknXatYdDxMiY6y9irzIoo5AuQtM/WysQHkNBpuYx581
7jAgK1oGIYx6wfjeD00xUKQBGlrzxohXa9dNaf98DFVjeKTDM5t64lnsbn1vCYcNts2ult3NEaiC
iWdyb4SsbAasbsYf2ZBsLzUuEm1ardQpb+YcksVKjlwVvzD6136ASNXZW4Szvn2yJb+hlhERyoPH
HleP8Gi8vcXQ5phPt9YI9IqRqUtII2idwak/id1ShERFeGHOYXbyrdWSZLC/35Do8gC003zUzSaG
grSlz4/82gvyPjnxFQMk8OBtLzr13ay2M7SSOwyF5ZYFxuAQrYS6L+QzyVsR+Eg7NvR1hpB+NyhX
elH5m65ZbYsZcXOQTgOGgyHsxiwLaCEchh+cPP2B5E6Qm4wodzk43K3Pt4i4qU1BUuWhsAKE4YeL
+AQxikrQ9BQ9CFQOeWiHrMGP3oY88PJk59iTNxw7VHD8NOFdUvOVcIn8TSSjp4UUtYKuIiA3iZxj
1vU90od76mLdFfFoj4Mj1Qajb4IfS81LNgNGFJzyDHEctCP9yZZ+OqwoKHRpvZygUCoiW3lS1nmv
J7eEl4AAxGSbH1c+Hhcb3EAimOfjcA/VPjfX3uLXLenWQtnsNCM/PMe+yTpEr3B+Lj0Cu3Otdg4I
coXzeKkyFEv9afc9HSXwKFUQzsU55z16AOES0QhuI0tsxaOy1ODj1QiZYMX62UvY0EpOs+e3pRms
9aJBQoLt6WsDJFXBlL2RWcRKOzC9ov1+TSiyxnaUlm20ZUL7quxSZKVQV7avBtsLAH9WWMOnTBxD
osNsFenjlCJnCdLkHZhjYMuNGIrqEBa4rMGtMMbHD9cQho4OI0+eMr3pYI0TzEfyD2wCICUZfWMd
OIYhSVXcsU3/MR5sAbR+KvgWfjBzrKVXodxQtFytzvRVNcWDU/EfpRY6y9SHU+vrCNEaRU1uJxAq
Hm6vJyxVmGnEOa7gDbEuI5PQm1PWVUvOX/ksrCQw2rw9aeeK1Q2U3G41DLXQI108DJ/tgIch94mf
jwrpd/FQmH1fhU82SSf0SH2AcRpVbhEiyOXUEJUFuIdKyIK5WXIzxuWfP4LRlyBJcy8t6q0w1aCC
AwQm1NpbAf6nn47SeuZvurgraolX14BRrp+nRBaLeAOGOZtp5GB4QbNGrGjQbGdd/lBHmVkz3f6b
6k7JFA1QgcOBkx8JtWON6i2TrxwwA8RlBBjcaBydObXh71qXaYSLl8S/fgclav/ok4rfGCcpYZqe
zR6aDUsgLRWmnimAD26jaM9PKoCD701/rQYXbwZfBcmUKHIpF/uHX2qeQztav5r8Tn4con8+3N5J
nliimoGELRajTyJYatG22ihYXua8TDmPt/bS60Ny/xEXdplS4oKGL6ODEcAUjhc4uKCb85B6zszZ
Lnn8twCjKL5jmId3qtGNDcpMA0EHsM4bycnxo6fsSncZjwqZF1A51tg3iojHYVruIIMOF/RDLdoJ
HgaAC5xGnyRRRktXUSnXlfwMdvTHCnRGJfKxCqzToCWZ+q8BQZGQEovBr/EVnYXoFhpGgSU23/9g
0Pqr0dYekYjo++n+7y3cgo0IdXEuuS0HOZk1eQDdI+kYQDFNpQcVqesX4HMgUrg7/OkrOfR4thSQ
KWy6Hc/NBmfdfqBpyPbbrUQ0fkMcBvvz+w28d+1y902mHuUikQYye3TzCUmhKmjTt5H3zhE8SG7C
HDVb5iRQ9ug253S7WxCVeBEiScNpOH7Oxkm42kz2jW8QAK30v7cxO6qAOLHPfjDF4A43pmlbpLU/
/cYfWFHZnZXo96AoMYg1YWMKCb7Gh5pGuMzL6TS7XO9BSBlDMatRcQJOOzNIRBqJqbE3GNOd1Ynn
5iPdbO8wc4PflN7ejOBkUJW6rJGR35/vtSqaIMe0GwoVA+y2KcgeO6vVanD6DL6bwNpaA8UepFi6
nNuXGP0Es6VlxC1gh+49ZkqB7GP23rP3WE7DfxSor6nbKQAN6UF3/55/HFOJhcTmLlkdCBBOVgck
aK5czl0DKK+h5t/ghm4++ZPoVTmjStRmh4NcjLHrJI2nxmgQAhIaB9RsI1lrJvMXo2gsC3AemSj6
gfPJ2srSjYEKa2fxUjncJDT6EeeQyH0RkxBMYFJmkOtRAb2+lxAH4Rn/8vVD+f8dBg38//bm9zgr
3zrC9VW6aVS6Eje+QpgGVjHMsjCCCEDpL6BGSWoHwxh11sQ0BlDIlJ269pBDora4pdFW5Hsj57Pj
hWqvxiOw2zQwKVZ+ItbwcC2RxD3px6kvMcMo1mzvaceT2A+8NB6X9IReY6tcHgjMbDjm36y+Kj4Z
VKpJFAMMh1f6aC/2Je33boai/keKKo+FuVpMcftQeis+RGZv3wE5M0z/jKZdWqwp3WfIFypqQQOk
miaummhrzUC7LATwA3ut0lEhKdV7tJO1hMliWnFS6H/LUvm7luCUSDMf5vPYpElB+IAlbAUuTM6S
YFr4S1Kk2Vhjo3BjpqMZ0TffyiWzLgnwIX2BfhpcPhlZNj6lorOnFNv+HrZySsOGk04yt8c/WR4k
fXtqfUrdk+6wX9jKtC2jOfKCTx00KQ2nT/Nii2Wmmei/ClBcaYLItPvUxhkPNQ0q66vWESlGFoQ7
JiJU6goXbQigKemEFStPpjWA34nYs6isc5eNyYArskVPa+E2/laRR92Q8QGpBQOIsszEZmGiEMtV
wrLxCLc3WZv6dl4PBshVJ6j7oOiKMGWlkK/QX3olZsI+3np3OUeQdnYR1XMbwKuFx4EF/vUuHmm2
ecQHIn2zr7PizUirzDEx1suvGb/dC9VFptuO3/+O+Sumb5rOwaQof2hBWmWCHpNj2d5s0zvnRpgK
fZA5ji7tp2kz5/gx1nGkYWR3uGsBVvyzSWCEMU0LtuxaFAfNtX9G7gegJgHeDSornNCO9Dj07Kdj
mf/MOcAQWuiP8VvxiHQThdnDik7uF7OdPnGpBggREqbt4B/G8GKG/14eRytwPQ3qtRFiqsXY2AUH
Ja36FAZUeDfL4SBHS2mHrw06tLuVUSd4eLzWqcAe0fZyfa9wX29mYwkArV5MFnnze8KzAvYKxhfq
Xnont2CNM3U+tkr4URr8QFgsl3u/eIKLVMuGAzHE8olSXtM/hvaeX88raylOx5+uCVlobGh7Z9Eu
N8QAbBDspddo2odn7grNhZygnU/GLpAFXdh5HIzfrpMouKdr6ieHJVO+Mnxklsu5A3LgY3jxguBh
HOtxVUFyEUZ55kK7aCBeyn1llVgflAtle7dBQTOvhN2DOrSnS9wREqG76p2hNp4IchIwpkI5L+Nf
Q+Rb/GMNanov6qhlkcnU9D4mcHXJR/Zq4D0173eo8Wn4VjvjX2nURJsXsCL8Qvj/2wnAZLy86qUN
mj0etr3CjWVjqEgcvbtlluzvdfND/WCMAV2sLNwoa4T/jD4CUvo8lIqEYEp5w+ElcJT3zAgAGzJN
TOJpxUD6yGq199GC0WOP4Xk/8PmrdSguFyAegol0gSI6OdP+DmCo2PzlOwmLCHbSuKFnYhm5L0+F
+QXrbqyv74hmICJVwIWyJUvYcFFGpsepifxNcw3Ua+vpfzqC68SMGLphJshGzkesGHiMgKytm+ra
3ArFld65BMyT/DZIHup4m+xR5xAWOEqPHDFdxpCKPfXre2Tfs+RBgH4rVqaGHFRjqS9TWaC04uS/
o71vDa+tRz/pLa0u8djxqnYPC/6Y2Z3qZ/OXegoPTmzSRUvPA64SVikYs7mW+d3qCUp43I1q4ps1
W//OhtKUm0PEEdHi3HWNW/V6CIri+kxoTletSjcE39L0FFR/UbKa3vNRzt+deP65frXBVqe9SwEG
Q85xESr4xI5o3yn3+uw0r4RSUdUBOrrx/PT+TXdJ43JcNeTMtQkONDVBoS1eUPbH25YMBut5chd3
qRdtClZoQLKPu+Ww0o/F1ejQAIUvMOtYLl6G2KGX6jI0Kjv02wzNwWw8QQ5lQe7sncDgmxPeiA33
8GK5Mt0rkwud/2pOpwuF7uEDXYT2EqRaBHGVYs4E+8OtCTYqvwdZ0AF+FzEp02paM+ISc2pMzlyF
mH+vBa5l3N/usBeFormisb5Stp7Ob9jU8y6kAtNIhG/wfa70PPAeMuojYs93Jd+JLgs4+xBRqVB2
cbbAPudFv8sKgjbl7Ppl/KXZSrOYvKSF8eLjNeLrsLtm3plixtTPqIYxmlM1Y0V0lAGjWfmxUBP2
1l9Rvo5QQLSsKdJqSTnDlqK90rT5u3MSmHYm5l+TZ759Mcz9bEh7zfIKwetKWGizlme9i+M+Qou3
6p6/fUft0J5Opgi30tqjHF8QaaSxva6vq9lVu+8LtBy2jSH+yj0kngVF2ZL+RPlikMGLkFGi8614
1DSupXTp5P+e7asadH7I4nwzrRVihvtVMT2Wk+iFN/oFb+Hjymllk1eF9ksuMJ1bhRfr9WDtrAVE
enToF4DnYuSlJD/w6n7UnU85TjhTuhfRrZNCHRGGoUJWYToDAczy6FKNAFGFnfS03P7eR5iD2c8M
9uhx06aJfQn0u0N+4zfMJaeuNNmdy+rd7FI+U+IwTxo6TUaGWNNarkL25+LhK44RIMVzgn55CQeA
SB24GVa6azqXZALlYwYbzRftKJHExz8vEAXSbZvc2CkQxJC7SGqYqWtnfuKiydRgsluBQhi6i5fF
5IMV4TdhqCJlVYXobRGTnJrB3StoBgTkLwe8uGKCvQdd2baVC5F2J7qyRwhVTQ66gXqhMldzTQes
QtSN/4cDWGLrw5l5SxZH+XwZO5+SKiorpj47Y7LYtypZDYTCxQSjX8ffSsLSwGbVf+e6rt1ueSGd
WLlV2rY0VYncKfbm1niW9dUEYSiZOYy3gGdLdQwyyWgXDof8cdsPTG9UvY3PvczMCnEZQYhCttyz
69J5WWFuJZycshPBoaRR/2DZX+JClXWj0vZH/69MJyEmupkn1RhynmGPfrGHxWUfoA9teu47XgUz
5/xcIoa8Uui+KNo0SKf7opG4wQBXaPuxG4s1ntUx6TX7s25Q1xY6+LtTN2xuv6DvGumfpgd7Yq+U
4kA84gZpKMTUMkaLIhOPsi4awrHu5uGuxEDHQsxhkI5CPhl1L1JefqmW45l8gWiTh8iRZOn8L3Wo
2zA6nmJogrVn/SBPi41Rce/EcRHJEXS3ZBuvg4/6fpJ3qzKa7jDxTU+5D37Liuzp6Ap5USuS+mAN
2KC2TvfVsLDRjzTrsNrFLUqv3DubBRzUSPV1+Rc1R+ql2z21xDcRcHB+CGhRbqinFkqqph+OxaN3
GeclkKmM2RANLWUhki9itjR0RpspS2VxQj12Ud7ldCrlnlQ9h/yPBcOo7ndS6c2me+8H64XBdczz
DFC3535RazcA4v5+OTbjZFO1uC2xFK8EL6+vKRK00GbMxUFyXd4nu7XgLZpdbrbnS0f/AmwS4ZJT
j3B6z4UlyKwP2y8eq2FesP/YNktUFVr21BLehM3ch7OE4gHqD4ygiY8eCFQNaAgnF1pinfE5FS9c
rWGi/S4oml1yGUmsgd93I6KBkcsQe1DvgxOODvUVIIrUfICzcvD26FyAmCYIf87FJHf41q9LyB7L
NUvIxTBYu4z9l8eDGb3XmSOh4Kq4xtSpm8WUxwGdhUyJpzCA4Pj1zObRl0+8u2zDys/PZRnViPK6
Cr1/QVLx/GLWtExlCAEvgLcdMLcjMFF+8G4/qTNFx3FvQ2K2wrYZBzmXIcFDgDbNJsYIcm1NpxBT
ylbwgTc7cgDnjodYSdM9LcsAvte4r4R9oDCL46UzfV4nqkCITlxV+nhsPCZdc06g+nNdz12UxLjp
kF79tTL5eC2zg3nlifgqnVWo8/uzM4E55pXvco2XIlG6a9rpJ7LFAxQUQuOBOeNh1VzvPX8/ZPwZ
YDXXUb5FhGUiMjRUoCL8nBLW2vQjRAuTRj7rXYOJZq0XFO+u8ScUZgThCUSvFpQAKPLjlQ/03pfH
aNiI7XLI76FmHcH+VE3DRFJyv/2kU+p+vTPtVzCl0LA0tj6LNce45HYQsC+SrVZvBnM2TNwMnzyv
MuKrzL86qics3tnCF4as7m5LatIFIR0qOPCiRf4FfWKtTq7DzufKNaiRP+085//YrsIHFiRoybpo
iT7ZUmyDX1UeXFsXzl8VcK014OLrvE7hxufZN33MHXc1Q9be3Uf7hgmHuiqxKCvtxVKC9438Homs
HBQHVkQTKErOHhPaycC/MFqeELPrYz9zzILajYBxjfQZjhPadp+nFIkeXR9zydaLxBr5mwGlsSQ3
lsE4lSjpDRnaqhqcaz/lVcmqmsApD1Vy/mgRP6w5kiE+IqaoXrNYHKl+WGiPCH9Ud7bfRrBH2LvK
oGiwQloPT1mnNN8N0TqgWR2LVZR3JxFaSlV1ib9hBDnazFkzOpC2/yXHgZs6p5LaQTZO0SmNueVA
NdSWvDnvTUztEPeIiUf0DPpKTbsrHGGD0MXq2kYWn9MMYO8qfqG56siwpRDWb2oTKnQOjaCUIAbp
ERAd6GoM52mLiMVvQW0Ey3xm3q0xfBLFlSC20SLm2TziOmtBwCZmgitPORQduPFIvDHmrJAbrOkh
fSDNqTc4GPCQskZL/ia9l34mB4VwgAiEJucB+9KNcQcZH1MaPXlDRWK7xXZ+NIBBZ0I6PcO7N/uh
/lPIqBVGs8rhqE72Fe+VHwfkamTch5oyzRhBozPNED/VzgoVMhf+Zx0VaQnA5UofxsPOOX5HbX3J
fMFbRSX8RJhyjzladhexTup7SJWwNpYYVDj3kEspJ4/eOd/oEMrReMV6nTEcnLdxO2P4U1UCZQgx
YF/3WeuWF06nZpPRnKTAr/WGbWL2diZEqD9W8wppO5OaZNNCdxQPEfaFWxHV5oK/dYhiPQ9jAUoR
+bAo8AtmVA44f8z73rABQI2/rDstKdg3ufnGmDtvnAZfz3A/ojMYnYQotJVvm/yzqOgovYYXwsPs
4V2X9jjgkBwiBZpf7duq8f2vRoOcNEPqIB/zPcZKXzWu4VI65ohfWm8DO29Y7P6sq/adSE5u5bLs
wOKBcX4NzNTR4U5p2OeWxLhOCycDsoQEbm+0jfBNcVwlwzufl4J9bq0TOaFR58ieHxSjin+RWTfu
nqb7tOiHytxgcUdO3YUivaZkJ/oBKHZkUw5Br0KezO4D1F4oRHntqr6Z9Uc/vrpOZ1n5SWzkuoNO
eE3JXa8fptIDt2W1zItfpFqPVLTN5MpXVkLB8wJEowJJPD1vjPdOkRKXVSKH06EwBuXOgvk2tJmz
uiSUWgXPJj85Fmj6v7uh3xwFYzPmY8vdL70FkurI9/c1eFcg4uyOUpyfHzmqraEDtlo4+ofjhDte
h5fpZOe/bHSxr00Pdqb+Lobxx1cLELxnGXPP9wMxRtZbDajFG9xha719GUGK7RHNABY/pAKzDP0T
bXk6hoYOpSiuIqgqNIFENF6hzBuFMPvIr64FKj9gUoXh5is7g22mhFvXcvlmtS+LRtXNHHSnbOj/
wn851ftXnEEyQnu51rlWuQdmDAM9zZ17oTdMDp+BVimJ2rhhVlduQ5HdLAXuEb4UyN6bLzAMMb+a
PSaFVegPKRHsNbzTLFDMvTgBDwiJuk6MQw+fdA05KofmgysVkEI1i0LDaNjsdD8Xkuz5SspT62z+
KfLzt0SVPs5aVPQAwDGpxThkOHGFE6J5j58Fu21+Xa6XpCb4e7blSAvnto979uyngW3kX6DJDeiN
7WvVq/eWI8bbGvfOjsaw3pWW1VZZAfC1/2TIX0rQhJYPoUBl3Qs+Ju9n/T4tUxfo1bRRMMV7QBi9
BA6IkQ6XlX6e39Wy8myV7dSJPja+uCkskEUJ5+FYOkL3XicIps2Yp9J/pG7eGsDeAMExaJYKFSbJ
JUpm79l5XlnmoHBZ/HPAVRmdSyYfX8PlVOFkyg8Z4TbQh+SFNZ5EL9qD+q/8mllyaAOFHoLg+xAi
zsuKmbfp5sBYGfG25nAlYmmeMYLVmQGAc4p/5Rpr95UrNDI9lXT+dncFAV8LcR4KY6HjBefZPTaA
tu4xV/sK+4tmGfnZSm/sk8tR740G4r510Oa+Tb5ErWVDnjf4SG1wV1ogimdf25epuyWocJ40m6SH
IG2ac9MhQhn+szVL3viNsDHdPsBVhzIh7dG4t62ym780iyPZHBHXU+Lvh/wXQU2YR/96vOJroQlO
SsZL/Xs69XNrMlMxrd3gTjqom+5A97LOsp7BKscSU8kh2CnHW26Vix8PYfzJ/KcqES8lXL4C7HOz
5TgMqOeHUWro2nDvEmrOnDcvND0iCdlY6egZFeHyIYZt8AoRL/Bl0NXkVZ8Zrk2Rrk8U4T9+ZEZY
oC2Dvsm8cnt2qwpJSei5RbeMHsHkn+OrdvcQPIUQs6dovhjaHSxSR13mF7/9u7KDYhY0WY7LYN0h
7GVp6r0/GcKSxB6w4HTw+f6bMlsnZx4hAE/QgpRMVyi8MCoUo+Pz331JGDy1CjN9igwEIaJ7b2HA
nf7HkOow9jMJa9jjAUCf6chSwxgbJrPDORXwb6TqDaKCzQiarGmLu3RPv3Ll1zrLVFFq+ctYvhnN
ac3L4cFVX49NdCx6g3E86mmzKxZ1qxbV5mlgcbs4ZmNGFangaUTi7+2PRmdSzdtllDvPWUDrY/70
SCtM5J3tUWt3LAvmjUSldXPz1vZhKxC227yuVSmD9kp1KGdE8Q4gBsl12lHv9JmcwnsG3E9sKIPq
dalK6mz2mi/gB7AY3CbeM68TeruUqyUZVwhrunhfVtVf3zJVIUO612dBwUwJAOotVwWcT9+4susE
HhYe7LmR4rl3BHTd1CNBTDR8hVT2moceV5btMrI7JbcBD98g9NiirzgvEnz9wHpUAHSHzncEMBPi
mHzQdft2I65j1UkSXwbKPeBu9zEzoqcRjkZMzxjojfr7HP/QpCFFj3oOl67fwWruxyBxucZxjjzx
06ysoCUSeNBZG+upbQrvQRTUhJIcLUIwn0OCdJdNxXwdB+zTb7yA+8bGGcpP5ruNFqHE4mcn5skR
kYfPhZNOm62MpFLok7Sz5gFKYzXH0JNBQhfUujoIO+pzFr8Ll3b8MvJT2OawSXVzGDONUOYMuDnY
mA0EXyYH7GYVMGaY2QNAi0S6hv5VPF3b5mqXK+u7zf2kdpHSxzowwy75mEDYIvJl8Id2uxJwjz2g
9GEP/6lH5Ks41WUd4uwuymg3hW2YxCRzu/ELSalcsT6YUS42iR0hnZJick1DdYJj5etX0sKT3iVk
UF1TyPKV3JRdYK1MHJifreTOkVZEW9/MaWt/3DmQhdKI8e8rsqAmJV4+F/n8XZX3AIcCIQhWqBnZ
vaBNcUhgT9vx3yC2yDvj1rb8OKL1veKPSZZeoTORrov82KitHnNvRkOHmEyzFtIyoF7VsgOhFSP4
r3BSao7L6T6tdLS5+SKjG8S8sgXLcqTrTODjuKZayGkbcVnKWoIj1DUkrWl5SMP+Lq+3Y7JS3u9s
zlk/+J/wgJj136V3+Ch9cYvQjggiopczEduW7jIU6LP0UqOqhio3SaI1HzANVKmdCz3V8VhGKhQy
IunCEj5XSWVutJNEnlIQecgx3bIOQkc9O0NxsVVCDVBUqe2nx+8Dk1cdW3JMnM6Ap8xLsxf/4NnN
1P/ZflsfFeDfzF0ODxOKcHy6mzOg4VAqMrPKBG/bAiE/JHTbJ5e3YUGnJ4jZZwa3AepRaSrcqnOd
eVAlL9ch+EjEadnymVejLK2oGpL7FY45GMIy12fLb29i7XDd/LNO1iBzFo4lY+eXwxNqTTOzrj8q
qi0Ve4H+JXJDtear0YgMsfKteyw4ORGUGL+1OBAg2ZeRnL4sUbjHAMplAkMsWEDw1zKET3aErLR3
6EDXh5u25VDTIsyizVov0xDlIzxhbEUkCuBVRREZ/B9rF3/G0ahT7AlH7QuAJlpdYoQykiNZL85H
9KHM2dbCF3j1YjnEXygdEVCp1XiB9dkfyO9KCmT/NI18m86OPXJ3lP4B/cIA+7wdoFTrGgnSGZDD
GLAJ2TeL+cdpfYBLOMtPLfJuQ3k4LNtmKoXFWcblqX/dZOan83CobwSafjgowX5Ppy2w3D0ho6XH
igObgEVYtCh/NTSrWTMZJryVzx52XKyludwidLuKlawUooZ3WYnOgUPy6cDKBf+tbVymY5WXMqpi
aJvEuSq2mUzTaYA+MxWdSx2IU+vBH5QkDsnQ/5tn8bAcmr59ve93gIAIfhbKeLbDIK8PXlaRGaXg
5piLHL+0ugbg5jfCY/THNGDZ8otAnDu9RGjyd0xSm0Xkr5DzQWVHmQyTUaDKQUWNdoJer/jTTGIH
NrB8TKpVrycb6Gkvz3VbnJrl+gUrp2StxUsvKoXhWb405MDQ3m79D5qbb1Rn5WulmBt2hZAoIMrZ
K70Pa75tXmXwrYpWYO5rCvL0g68Ph/Nb2+qz2xp4f3QsIDt47j0i2m0pRbCxlVqVrWyllvXmIGPH
cVotYKi+C1w0FwNg3ocTD/m4b+REeGvVMGq4Hvjjzn0m2ziijMEdfhWxN5LtL/9iGLXZWVygrNd5
g0yTTrc9DEyA38vnPTR08tDOLdH+Ko654rWl9NsfspZMR5LiqUso0e6Vm2N05TadwoWsUO7k4FWX
olq5YTaET+neBsTs8f5s11iwYEZjmdN94/1Dk4SiYNXqoRBspqLJNe5TUSxTwiN9R0roRbiBhy5V
U4/xUPi1+eGjIjK7L+3w/FCmHmApQN3kyW/pl2bl1gq8o8YFTBMLwrbhxCWjIx5dJKthR++vEUSw
DXMo9gJK1ldRVSnOwzQvhI62QQokuWWEK8ee4AjLfLAFBPnCPRyvUDDPsFWe+HM6/x1blJwiByQU
wXS3o9AFMHvfw5XSvM73gtSfRgqxXwiwRzKa+nmw/eY4mWno4LwVxskcOqUGJlz6gYmCT4dczYEO
u053FkU25wqrpx60RFCTAepBbF8M7AUu1wqHSLp7r9Up2gZs9GO8Vlty9QgTuHgjFI6stGK6oKV4
1cIcFJuS7xsmqcT3uRVKxx9k1XDxYieZyyGmoumU91ttFC5WO8q6xOhwwYdrgh3wc1vtSNsLqfGR
GDN8kLmxx0kIHKfpuEbOHyJCQE/fH56U4vCSvDoDM8BsJdJfvfUE3ql6e58Vp1x5NwDKS47oo4bY
uNdPBKFXYxgrwP2orhOVLcBcp8brlGQjlNnDT1/QPPC9Rvp+e6IJWayooxfysgQU3NGbAysMO1mg
hnxMKOmrS65+O3i9ATr1LMnr4zBtRf4DhMUhPOWU5DyGO8IdhGCYESDZkWDg5ABKnMVbgp+YWZa3
nNb7asoMyobH1P/UY7DoUVWEvLoPx6mC3pW6vnLWaxY8uniCJV6NbF6kvoEJvOncenu8SDw+PXFz
iGX0XA0IxRKggEro8HuP4z7A4/AIe6UQDAdvUYVT3rXVQTMe8nNZoGtUP5E89ofNu3ylf+0EkCna
0YPDvhYjellAUXLwzBrBhMWevRNoQVTZdJ9//svGDPuacPtpbNeOl+aemivQcYjNVe50mBi6v7a8
3mR1LXCS2f4CCCZvA8HZK26UYfP0aiw4WWWBXqMvQpNcydkzp72KQnJsYV8RFATl2XsU+UsBRkWg
r6xeG3/A4Jpq/GMmLZU5/THpT3RxG0wtcQ0SfI39Z0euvknP98MoVdqTmeSnmellGPG7iR2w4tXL
qV+nm5sbNN/uF2T5hSj+1hx59F/tZ81Bc00XVI6RIMDGSmxha7MuNIeImK8JtNyItdYcWyhm3y07
7Y1sLK3dsrwipwzplg7ZhAUAq/6QHnjwMqxtP3OKgWV3O9YCAWatyqVibi8OGIahIU5d/lS9qSaa
yqH21j0vgF51//EvOZRSMeEI0euw+geDLXzkrMn8+N0xmjpn+W404sxRsaf2FAEJeql6LV04H+lU
0PPowW91CjiwrOX1EWn/8lanpM1fanrk157ZY5ggO37c9GQh2eXRnFiJk7HqFQqvVR8gN+fk4ULA
jzBgj7pQrf7ohCMGRGJOWivADYPjqC74OsW0jasKYPYi+pS1xEEKRtg4dAR0J1pVCqyhxd4EbZwb
ml0C0Q/eQksXAKxoizVGne8jBKoC0cETKzYJmVQxBJqXgDY2fB4A4th1uDaXxAvll0JjUUU5V+sP
LOdNn3RAsnlLtibu/V9I5hWuMKbe/k1BQWJ52kP0yaFplcHdsDFurZwJBeYMoJuOsNXXQEh+Y5ju
fAOuxW2xggCd4hiP5LvZPkXRN1U5+nsKr4VVl9uvv5DZRQntjDkMIbS6UPV44hREetDP8y58pAk/
tDiqC1DeovqEDF2oB/LIao7rEb0BsIz1cMS1w5p3h4K6d1ciYOai1JYbmex7CZIhabKC2b7bSXHF
K3HkNrAx+bBDnprb/Dru0bYxylkIB49bzLyzmlxTM9vE2kXBMpI3DjOETB0Z2RyX3NwZr9BNZEwr
foszNbw+LaALu7IteuIdeI1tMgib5q5fnKV5f0JNev49sC9Y+17Y3npRgywVVEwzzL0z1P3z7Rcp
WzcXF/lmme8K7FtnNX4OAAadSi+oFbTphbgZYV9PfbEmyb5UDvByyx2EyCYO6xLukKSThE7yUSN0
mk5e44r43ewe5VTNY4Rc8kAplS0l6/+DyC9PoZCk1dRuozlb2wzqDsFx/Vtd0uvJzweOk0XeUNLz
ZQLGD9IQH6P+IkHeDm8ls2Ef09FN4CfLBkrIyYeKHqPKjNkfA6FcpWWEmz0EnM1LfMC7Ie16LdA4
KCazQxsLBXiwKkjyejWvnY5oSPNQTCxS3AWlx1PqFRuFLEY4pVsX+EJVFmIOZYliSzWrVglG0ZeY
dRQ5ct8nuxAd8AFMJiZaTovu8TyDhMIt45XtqBMNmiIoe7huJM7RvToFXIxuNj8nsAjpD1Fg8qZz
d1+wcVYQO0eGCr99nmNEwctzoa+6fj0JGshUvloseUbCm4LBC9D2CR691cDmtwp68+2a/2IW2+z0
3sutGruz9aH5h75sL4yUQuWVq+/z2QDNAzcOTB4vnEFDHUmwXDK9A5wRWuZUD0UQsUc32dSyd6cN
dP+qoJM6of/v2RpNk5gjA56j2YDELxp/yUyfHjWKdG6BsW3DQLjgmISZZ7uUVWCUF1IVfObty1+E
qCfsvMgo0fg8kxlzxSeE1C6rIsCa6+XOtRKkYGd7pHwgEJE7AzGueHoavHSM+vlz/9a9kWDVX2iA
LzhBReX1OzZrcMQzvhrc9bnWt7+pi360uKDA5n6wkoxN6lfxMS1+IKDiBRAIloIqXSSYjJDgnp+z
v0aWjxRov+dPavPyJDlilIVUA/hDYF8vmxZ09ueuiLMn+rK+o/zuP3AoCS49UpyjkyT5iHG+fKLL
FHET4ree7Ed4awzl2n+Zxn8vcwJJ6r1ZmqpZ6EZrKN4/VL+QjcU68VuB6/zH5IGTOBufcHUy41W2
f7M8Mdd/hPvLPFkeXp8LsJB6fXaIuPOSVHWhMACbHYLowd/Zmw5QvPa92W63RK4HEvwjvzaW9YNe
74j38NcACQ4VgVKbhMqMuGPMaoy0Q5XaaCfAYEZRmQ0ZhUXktIt+my3ewbuysNX//01Sulg/CUGg
1lBXTMziDERZALsG9rcOCGSBExU8p8IjqCiBoVKdQXfGbM+NNJShQeWUgOuDP2i6pY+wCjFWdlk/
9DOoKS8Xrs8Y4HptCohu7DQj/4bcKAgKqBooTdxp5yti6cMt8y75syB/mAF/Oem0RHfy4XjTmEaA
umAoza0ONLdkr8fdfOmVTcRL0v3ltZrTMD7TB+tCyy7qM5FA1BQN8leVvihTMVniv4IMfJBl2n/C
jpGVnFG7czfG1o7Yh7cMBVYiYl1cfobgAGM59W1PfgBN8h8dZTELUrS48qfgo9lz+NO9GUDKleXK
QAi69fEVXUZOP+hPq3yK4lNWya7KH16kMUUpfhJ19h8ED7LX0nxA146O6hjIU5BZg/+ee96O/kZB
397xLMBYWUa5PW71J9xvfzIxIOHCPvcWFMJ3Ur9rMPvaUz/qOKroYb9uVmzz13Y3KRsHHJYQ75ER
mejQYV0fPN2NWaUJbQxerKAKP9Bi0Q3WC1dheGX22Ix6eVOqmwrmpCPNjQU1ZWmlRm1g1yPmfqdQ
JLSsiyht1J/8opI8D/XyXfyQ+QFxuFN/C+cFTdCs4V10Qkv4RbuU3F5Qjlu37edmVbyjGreRl/8L
rGP+wdA8RnynHOZjBXwdaw9FPHP1SVQul2v1o3flVd26fu/rLxfDDsFtjiVMIZXZSa5Qc8WIjCdW
/gMDHDwxQ0gqRaZyIOlsexH1JAyo8avjFfPif8mSh+x5r0vZnATyBWd7ryH/cipJq9YNYSnWv8ZB
wWMKPlqtgZVKsYDwM8xABP7+o8EsR+5cU1vtAId9CWmWoZYcs8Bdi9Mb064QBdhM5Ocl3sGuzoEJ
lsfBrmpq+E041w7oSZkYZt7nOxDB/ubcj8oE7gQJL3zVKSN9ghTk2A9qlrYq9MCl5JQKdrVwGUjM
4eCV8y9o+6BijZlJ2F3UTn1nnoN+uZiRIiIH+oFOiFmxkZdtWbyfHFzlq/Z130gFXuDyLTM1Zb6K
CthiAqls0UcncAROomI56ksh/+5QzeUQM5wFD6etIDwD57eOTjQwR1JpKREi7YF80eAUfH1mBG/E
ILWncw2xr253zKn70R+W4a1vohLCEsuGUGBpWR9ccEl0OyqfYnVpJ7GHG+dY4OnBGK/lywdZ3UFo
lOn5I4yxxU2qLZLar/qeLa/yXN7pqcVIX5MYsdk3dY4DTZvrhQRJd9LtMdI0fDolIjhZUaN3mwjF
qXcejPnYq1G7IuV29g4c4N31v+gapkinyHM39mIRSo9FU5cPVLwqasNVoSCIseWpebx9R1Z9Zu1D
lL49Ssk3ZxSILakrNl7dwpi+FQf+tRuBmKrV+mnQLziJvuqILI3irYhLq4DgMEO6ZYEKO1BbXnE3
gPZHMWGSR6D5Qb6oSYq1Hu/z2YJ75z3bqhF4PnjjYb8hn1qShEuk9en3Q6ygwOxx/0RfP59Ls4te
F/XimcL0ifiEA2A+UUMQbvXkdmBMpVN26aO3oUrWJSRGfc/HIqXIuVW9cVEWJcqJHckhQfIaiHIu
2vOMlICw6B2JYyRLLxks0XI+mQxURvWnNho1NiaId/4akWMtWXrrUqwaXDssMWPOg8csnyNYnkdQ
+9knyZmT9RwHB9Jw/cTZu+1kVMI1ZhozxjvRBn3xbfhsX0iFFvN0XqkAX/xusPGW4qGTzPtacKR/
g0QS0MOGpnfKS0IeaPrY9KRN+88KpS7rP1QRifaqHEtldgb4eigrDUXVv0N6Ns1ELafdORaTDZGa
LSnRW59aDDbTp7qadv3/neZ/Bvf7dR+GFysNnAxpZeL+bytlETt9U4USns+rmzTfSu+HJxlyZuaE
XbRIQ1ERAWuBISUHIEkth/1yqNYN4BDZR/f9QbxvdfAcknS2E4frF8pMHBnzyuYWSbEB4aodIm8w
y3slIetelXJgYxMEPJAcOi2z3iCX/Fts1l7haAlA8MqFvYsqdbiaakAS53fCHu1glWt7qW85Xio8
KtWqaYVSmFtjxOQPNPpcXGFG1yQ+4fV/BqNuK2oKzcap+Au6HfyV8gENtRemGiQ+s1AzdupiBwoN
WxFgggxHleechq4CuqMhdwqLEPz2tGkP0BSG1JHM0LNnF26I3Z5wXfC2IAW+WW59PEMuoDFI2GZv
AxupNbVqzYb4q+M+DJ523e+TIHOAuYLDw83sqARk4mX0hNnAbpQfZhfXiLd3TXJZlBJkVFF4wsL2
Gh2lSPFko5nSHRccpPG1IAW1rGehk1VCsLETlOam1K6XmVPWzhopfUXyCu3ReDlrBOD+c1e2K5Bj
mXHtlYqkNd5JA9v75uvOTto96+SU+aRK/0Gl6qWJmRSIMB0o1pMuRYC1+AawfiLbt1P+LEU9dqAB
Ty0640J5MpLXGtmaTLR4m5qMSPbJQd/gh8Y+dQxrlLko6S8xE3z5oNBHeud6f1DTQK7cWX3kzWdO
wVnALC2JTCwQD+IF98jjM6qVGr5pOpp7/k+UyM4tziDUOg1w7gYhzawRQZE1Lu1wA3jF4pBs8GlA
EAFmuyzPLpfvTs0c/iZQUH4Tt4QO+e6HkZzSekrQF6ZoavrzY1Odn2e4LYg2yE1jTt/yz4Dou5pA
fcgsD/ARn/3D2dSfvHBKwc/IOu7uwNDshCVecWeX/ocYO4PWcJWbKJkGUoTR2m/1vq4WImdqHenS
u9oQxcNGNs6Ha+qsH1lTr1TdqqtzUr/dNRxa6R6s3TgPc/pCirBleAayAXL0WtCooufEXiIas1eS
nFxolfX+JlreOmMe6EH8qndIKUs3ClyLmqCPOg2C+sfTDnCFx8ufFElYRSwQ/2MdV5pN1K9NAuIg
aO77OTlK3AXk1DQoBzTWJIYFos5WmeRRYnIakhIgGZ+eLrk+mUkwMud3PfKIgDL8XsrSbBlyBiaN
704J7F8JMnoW2DDWbDzrxT777DIOfS1NHK3OsNeL1RvHl0KiRr9IbxNo/A4KJdNppKOhCGb12K2L
5KAN8MfYV/aPeQzkyYuKHm+hl/rcWGqg77jltRGL69dztfzOwJgzGDh2QnA7MA7XKZ56XR+Vv23I
2LFG3//D/3aVNuz4JFzUZ/D5tJRLQ4RTfTYmVIHkIiFdzaDczWoTJiMxQhq6XPQxZKT3uQJlZMPb
LC/hCQOFjM3BSQ6iMvOOkSVwLcch4QB+LWtFyRAfUf8+OXOyrXWgWyjoYIvcbN21sQ5Ys07Mvp/x
33GIg/JfaIl6b2hTsstVNkd5two1uJaYFK3EfngWIBYLnbshRWsTW6HJ/KH4DFROmN/K9wLm67+R
eDOlJO2WkKnoLuZ5krtl+fw2wE6Hqk/wE5mf4K8onKTCutca/KckkO372zg7nPW3rmfBu5kclbgA
/kGDeqnLqQD3Vxucd46TTUffkhKQaDujEFfZnBqaLmHqWJK9D9mhnfHXVz9LourvcwVMS4Qs4Xb8
Yq1Pnzy6XWf3DzqYEOUQxPPHB9ueF9NGkQAUV+Z/ELrccEOalhvyjf/gdzSg3VaXcUrVvRyWDWhx
wRvMvEBw9hKh7EcCyzSOGm12I/rXIZhVMjmYdkrpdZAW705JX3mrC0n09Xpu/gDxAoR9VvyHcl1N
BAGQ8gsv51EoJBCiPLN4sOGS0UQUb+doEsj5aEPwyhhvZe+1d2MWFRtB8S1CMLiCTdoISy4oE2Ix
gKaHetDb5lz4lZn5fyXFhqlJTxMaQj5GshPP3B1eQG5tafLeg/AQJMwJjqgaczlfkbM+XJCCQJNV
a4n/g1wVskGzRj0SDm7hw/aml4oKQahSEX2U5KYTO6iUdbjjlYTNnJOzCbkjhoTERvas2zbf9c3A
eG1+QUTpl+0LSavw7ylYQj7ywzkrTv0AZscnFAiqUmROPnwkD0nRvK8WBY6NjZvlP9boqEIvEgmC
MrJPkBjssx9yuGIz5vi2GfewmfaD0OZsfKBCbTkqVOL6wGtUg7JrmgaVsQmgbeWjy/8P97OqU/eY
YtnsHcPTrJeym+lqx58uGaWL8gKUlIl4pg0J7asCNqZCPL8jG/YE+xnpAFnm6lN2e3AqvpVilcHe
k6/EDxjrKftPYRG/x1D5uBocubutmcvNFsUwrVBZ0YABXhmMxmeMKeaMONDQwoh0+QXP/gPcwiXo
OFEFIr8BgrM2O9rocZ4wH1FI/DU6yRuGwAbHHJnwBMZUXYrnefhW/F65+RfnJeuHu1dawt2RTQ5E
eqIv4iph+1kgvLfkDVWWCiOjKwiiAsAoOWPuXCtzcw5YBbfTQWOI6SbhDcDazCFFhlYY6N/K/SHw
IfoX6KWYYC/4Zr0XJzXae337s/EY/n6dCgTpF6re5aSAkTIsOUzUrtb3Aj6mmlsk6yUyfoS8BK6c
oML+SJJfpKDxuQWveNAj6TZvuq+Gruiiw9M03hLzIj+cvl3SwgSsxlzUV0dbSz16QHpW5jz/OMQu
MuZLIBeEkUsN2Bp65fI1YXW7jAZZY/uBN2ZqkwHLqk8UQ7Tcc1t9WnJ5ZY9RhKfkAzY6wWCw1fNY
3lARFk0oRGp9CXLr2w+7ClyUnU0sRKEUjAf2Lx0eV1GCrKEf/FjHeWyH9ZFrFaJKjQabEy2rGoYe
l5do3mJOPbj3s6wF4qPXwWHfavd0HPL20zsMJSc25TSRv04NDmHarZaSwRoNjohQ6qKt1nXaswNe
+/1EpB9lZDl6V0AMd4ZcE4YPNtuAxp/IsxwHKyBOWUdUwZtd14e9JLuhhVyhvAWvAMP9AJhJMU/m
4PHDeUvM8bdbovyGS92p+xUUQCpAd0BnnmvsIAE8k/61BEyA+XvHT8hM9XkWkmecAPzE6NWzxNwK
Ea9rh+kE8n0q6pqQhcre/6KDE/Lv1h61oVfY1tuput+ogZNYNj4FXClfYN/jskbLflVYGdPs1lBw
SWPX/3nWJgB4EqsjiEKw/sN243Dz9VLihIol33sXsELjL/1aaiSF004s5tdKUCsVUetxdUDgkY7b
E907RiCreGDZs8V82BW/TMG2GzUuao0p9nJosw70p+ID5Uev7TrvlGv6XSG0lv0Wr3xTGWFNFRHL
7HmZ7N1LnYvjFOUmWYvIqAq3RVekGV02Rfnd4v8kWV8cWAfA/jwxBq8exuoumISo6SxGzhaX94pv
k6yBgExK5vDwxkGsnkmDG6oJEC9ZqW64uO7AZla9F+/cx0hujdEcGn0IJxyMpqRM4byAjmh9ClvQ
W1faqyZTqMAWfjgJA/vgItYi5wO+21p+TtIV4NcxRLf6OJoczar6WpR6GrOrjl9BWzTe4jYuT415
mxjNWetw7ZU0bDwvAgBmUwb7R7x+2fJedAs8wIAojShy5+BgznVq2MXAIAzhW1SXIv6e9LrPKepL
Pko9gDBaVC8f0npuQ6hcKgHOm9K7w+ePf/hx/MjnWWt91B4fBWP90/kcBJ5S6AeHl/emkrcE5rp5
RDaT3cYOS6+CJIn2zcku8yMAt4LNZIXmG1ZuKw2XnTNi3XF2Xur0UYk8SbW2EQchJIu60B7QA2By
5kmJmj4+BNUIohrt7bKTn9gDH8t6VfPY5mTkT03a7Szs9SRnxF/9CjEBi5C7wzpVb3S21EvweyLf
bVlyqPIP+R032cEq03mkaD3mpEv6/ZQ3IuzdHQWCTgW5Gim/1bIRxJ89ZhmFEdfrMd+lSBqzGZK0
pBeMfdJmLJu0ztIfpaJ1vwH+QjUVnhD6zh8kUuFkZ35xctA0blMkkDFmltl0As0g8TxbGGZfCQle
mAac/X9HoG/LrcILhWPeQZ/S5tmmj1qfWWxBfj9WgNQMDGSxoF7szwcBRDYX23ijDVakyWXn4ap/
zZ7ixv22sO5m2GlT1kUoZJO0IXoZ3zJ76WtVs+NdrMySCWuLQAmj7V9iKkgTULgF99B2zbqqZ6uR
1X8Mkpg55bfglR2v+qhffj9C2riJc9+WlsmzYq9qw+jx/2hFUpT/qh37YXs1yr6U3EZ/D+rlSEoU
v6y+tpeaQYxDqQM/L2jmL99EdEzKP1zCvSTlH3vD8kHD6s/jqtqcun5qk8XZN/Zsms2kjGqbrIXl
1IV0k+/YZhEVrzJHufPvNoWKkKQyj4fgNoqxYG35D6YZ/BNWIEEPKOxPbimTvyb0iRBCek2PZ8xl
vfUFNJJQZ8HCNxepIhrqREriGvP5hvHeomjMr9Yy/xzOqCyyVd+2j1QKNipOldse/VZTd5pglzid
nm8kmn0sOAe5QRing/bcMDCneaLJqI22ywNX7ogjVVR9HppNnoMeH/vuz4RJh1CtQHzJHvQiiJTn
ctL4M8KKw7CtiQBGNutdwA4ELHyQW7/PzPgc9/RBteD2E93+m6ndT3yZJjSQCvsc76rq93CSkolY
c9GObttzGNzDlqePJTFvtKJvQjAxuo1eCCKdkaxDa/H7uG4A1QkIVqh645yWuRQ5+ZmSj3e5zNNg
WLVPlvfbN9YR1n2g6wQSQNWiUfVxmPlrxMaG7/fxF9BUYy61lh2nWQ1yLZx1TLdVuUwLmMupoyD0
6se1YHlRIGHb6aXH7KUnQZO/QUOylaBuK7RR+xXRTLi3xbAe92/zLwPy3/9JAUhoP2/BZQtVFkKa
Q8sjfhgsPh8xlhu/DbNibjuvWzQQHRlrwQM/XCfGqP7TBkf66aYMfyqQVrqGP2m/e9eRKbfVErd7
lvKYIa3x0AVtLhIt8qRcd1kU/zxqJSxLOlDAttG3JdbMFEk++66tDrlMIWwzYYWnZr5Wy2n2rHPo
0XzsadODzzd1HOwXj+3uHVUHHF+MfHZVJfd93wNEjXlGKMUtmpx3CLsI2YICFvOFN0n4XGmRXT+4
Zv/KiU76abGLKUv9qewXnMThF/Yag4IU8zOlaNf/Jgm9QgfUv16Q5WFGoHNbsxhW2EIkQM/7xcr+
5dAKXr8FlF18CWJnoyKwNbyEtZkBonFgw3eN/UhQRFLdmUSD96YPa4kmYVIJTYvckg1L+OgXdc1J
B7x+DO+GCTNTuy2Tg1/QYHMhBkH1uG1lEBXQcqRJ4ZhW/xo7wKC48MJXEmG0cSQPq5b+l+j1aeNN
BdJfkwOkjs0XDTdRQcVgW+5E5jC50Cinlnpp7yg2/VRC1/LZXCo6lQ1fHx9jga62nUwZrQsj+gd3
ywmEiX8MsFFRMHlWa7mbEMkrySr4y4Dmdj2rAdnKyz+8qZUNiWy/9ThasEWf7vEcK4H13w3QCpa7
+JYflfGzWt2IG8U2mIS/sosPWKd9AxhSF4NM99e+bCN1XbgaKJta1IEcbevD42NRMu9d+PQEfKJ0
nK2A6V1I5nXuMLJ+5SqbYp9bBWyVWOJVXBTapYGkQcBXIThfOpQURHzWx8jy1VN5el5XGzGUfW+D
rpKDyZiPTsfmSv0VsbyjiQo/GEQmZcL2/yFo76UwkoNn+lmeqf063S/AGSf/4NdtE3sDit5Uhj9v
8MhDrPr8EuaYR8/H+Z9oKOgVty9akeya7BSqDTYDtTFMgpCpz7210kl4fIfuWgGg9SgabdV6lyL2
wG5ITRU6I7l6gKOnX6uQAMIj21N88yy4yrTqq9/7rloT1z1dCnZC+WjqvK2ZcffDMWGgQcmpGTM5
42z6NrDhOeSJvi+UiCOYp+YdBzbDLvA5wtQVQGAjDABShpCTKIatEhAoet/GY1hl8fMiCw773lQo
HPNCDwbOPc+LHqoOOxUWJ+ivvW4/QqyLA/GctK809ZWRzPLgD3+FqPByyXDgmPEI3vhVJOgFL/ig
fffaTMI51wNnsLupQmJqCSR4BfkjEOVZ7tByOli6lCxkLMvH0N9EjzLiFJtRMW/W3SjIZiwm7p+M
HCNF6Vk/7H4yelBrSWctb+JMWMRL49awPAfaClAlTuHGp05y57B3iCah2Xiq9sobxKeTV1RCGH7Y
f5sy+4HKSJjzwtQvn4TzMaid+mYwvNvuaoszYYXN9ridA2nGKMOAx6IYuTrDMC0WYNCZb4lAQ9cH
kRtxMjjvOx5sLxGEDaN7CYImqx3vSH7rTjUXQRGdfLmNij2fVpxOFHJU5CRIzy7Cs0qeyRdtsAHs
20wJwXTrHboZQxyyUM7HXpvA/SdYEnVYvEbDstTg5V3ateBI8bH/NzpYDWXPcYkS1gN0o8RmEqE0
w1h+tJs0+7uKCBkOYQC8a+7ZxEYxxTx1HkxK3UKzcHLGdRiZC8bX210EIi4QjZ0hTaKXgxlKPHhC
YCcQmIS4UxywSw0DSqXmjlQPBK2zz8mdJgM9OJ6NSQ9jao7u+ei20bThtOt0PY/f2mvOMr44XyCh
JENQ2h6jq5+b14N4erc4U+aA9xYIW2at+eX6e7SmnHmwkA5TW3wvmhNOaD342MQYmKXstR1udyZ4
VSddQA1tQjGaFP0qc7LeP9hanJg1JaJEQcg3dyhxKCQ9dlT+3RJEKL/29xVFd7vqTAFmsa8OktEf
z/+MpjtjV5hcKSaAY/Gauvjqs5FODf7YgpfzyZrlvHJc2izESrEbuvyxfJgj6M51183SmTVyht3i
qG/etxJ9iRL8f3wxSaF2R8AjpoId8QXoG2nniFbk7pmxgTkGGbhli2YPJ8wYn7LnN9cJmHZyEoV2
oIvo8yNHQa+iBM7VZUJxxCQVU+dQ2B085wRDOu3kXNLXPuoBFZZ3b9+fgLtuIG3qbT8ZNSIgUqDP
0zJt3/+mDHmbS62CzB4To5L0u3jWOysy7ZdkUlBtglZJmTrIy10JqeDC88Tm8grqQG75NCra1nFB
czV3LEiHVC5ZP+MVwKu4c8m9TGDiAsMkuk3pXTdwRvAL1FRzwXRoR4ctH4IbkKFBz8OBBdhqSPm1
qNEfQ66dmECNjDXL4pMf7r0CqsuNSDpLRkPiz1quwEsNfvuSBTzRNJmnMQQemUoIdkOjV6jqwbfL
a52Ioc58Mmv+sWSISAyIBcoS/fSVm/px94S0jwUdQ5NpClpZ7eBx0qBj36vRAK/BftTjxc/xr3t2
L1KjSZDzBVgilEwrWkY13oijl3xL4+gtUKvmpKot+b4g35yHHglJ69ds2JHSkSo3FAH3PwfMuWdC
dNlqnYRhaJYtJrobVZGGmNNAQgeIl6mgy/jKRlj+rjy8q4t2qrqbjozMtkUDtuHArTDMecvylB3X
Me8cDSemEM8fFVzwZd/G43Dcdw7see/JH6y+UaWrDVzalqWfmr6FtqAY6jv4gaTbQQKTEjXRBayv
7kkMuweQp9uG/MBPpVnRhoCTG9dUHhCropHpx2LMwEhtCbfsCclRoAoHj3ZykBQ3LO04hjCFIYtW
W19UXh8yv2Rem3ZvL9/g/t4IHtdQskKnrosHEMXnq8Z6aqSbaVp2VViBwQwsh0jsbWzWt1W4RqNh
l5V6K52eKemd5q/65PW6c2oY7De86OQQ9wVWX5GWtbaAa+KLdrR5WewO2ka8JjjBq6tJpQu3H47F
FaKBvNMIYY6Uk/kx8naSa8WHbCH1Uev6QQY3FRAgqLegvzR5JyUiCVsk2RKTYUMhCy4cdQJ0GL3b
64YtVNkSas7In7CComns5wCunr8FDlp2q6bmaiKi3/h+c4bgWJWxt2g79uy/kQaifQk3a112tA9z
L0ekVSU4cGhLn122D37g3MOX2xto+/C738nzuzWcSb0WslmDJrioNi0gRoi8AjI4Gr/+4p90bax/
JI3LYcV0sNkkjjLhkV59IPtDdBC4ngH8nEnP5UvI3tAP+XOSXUKmKcPi874dXRSgJmPOQzAETmSQ
jcr0MfCSUZFJ6kNOe5fb7MEpnrvhyzZLVZ+qrPGcLPRk3kujF7bgWDDHhYV+JuS63airbZYry4xy
Ac0BJdJm6CTUO23nadQZfPvfJWzrqsu1vhve2//gAaiTLY8gk0vnmHvkVpkIYPht0u/JgKjVLVdq
DfQmwe+RttlZ9R/auWS3YvhgeNL4xdus5e00V0cIaVXDS6P3RIaNBEOvluG2fhDT3GnDNWaKUDVY
iL6EgK3b4BEknGmJpLnN8A/fiSG5iXj+U8jky+kxFiqwRPS67YIcqwucpNsMkA3Bav4ddwLdsvm6
pqYjppHlIqxcTroxTGh73TuaspxVfNXLFHGU9+sTzUtKdRNodb9i8ciwymEzzQfvKuVis/oOs7fo
iGBnStXGH2aMhyZYOeOMvK1iWqIyyP7NIgkmgxZZM4jmP5Lh2BT0PYwc9U6v3I8Cw9scArG4Ijar
Bp/RdovGGXvcsuAH/laYXX1HniQl+AlE4ouEleqmp5WrUuXohQHqLOWZY8yeRbfyfSfART12gdCM
4KveOn317nsiKL3HJW0z+NWaca50g9OuYmB4H353CPhnTIkNsRUl611+O6BJrixdtdCeCO0VmzHK
z9rHXOPttj5RnL+JUVPuAEdFMoKlPTvDV02oU/nSNwLRVuQOz6hynxh2jPwVtC5LcBbLeZJU8dLy
FfcIKR3xLdpyy5C9nrRop9SE+1iSbtinWtJ5cqCBebAW5wl37D2xQwJ2tjV+qv7h0daStL6Eq6dW
wpvQWvNmZ/dEZp68uoIODDMYxmF1MM+EIjpsCEM+VPtrFnqTWklm7+XlukTrLIB6wJ6rjn+DuQaM
OSozVA2pqOuCeZ9042cXbQrcVFUI318Yn/RmYQ0P1qzJ9STvfUFm+apxztbxoCratrwThRkg0ZzR
h2pGToJ43VrjBXCwgArwCJe4krdArVxfiP/MLapZuWmzcXell2xYcZqQoW7XIXbeyhRLjE0UCGxY
MoPON2zFBnfBJ630xDus0LKF6rHGYu2y0JuauXDeXn70G8wIBrGVusgckKj6WjuCWeCnRuwYy7Jb
gZvqjt7LF1CsPBtcXMBVhHZYNWcYFmd0+ROj37p+55/30OGreGg3Lbx/ZHm+uf88MUZMljsbxu4l
10kxEAi5AJbGyz8skIt0xvsBUd/LA6K4DVvnp8StXemPkKmEzDg0Tg7Q7eD+YU5i4FiYvxht6Gjr
R02g37NrYxvoyAVIQJsBVMMCvIef6Ko18BDSCZKQETG9cgAuMM8m0SIvmutS2o/ZVEDtLQla0WIS
ApNeyNiOoTieuziOqxwMGNv98S4rhegTt7FlOJPkUChkz5ZTokdv2Cb6P7yPyjGT2sF3RflpQmjg
+ZNmEcxyHflM+ySEIG28AlDBkfMt11x/Rg4tJDGytIf9NNWW1QbPfFOjJVTNr+AT5sbLT8IOpoVS
hgKq0SQPWp105NZkSbNrMeVTor/1efHJzgZCCY/wr5K7RLa1tunGvx/Dd6W1VqRBa4oNN4QobtWl
EapFXgvzk7Lz2SVTRQYqTW8UfbSMVqoZvvtr1SJXBgtWxj2l0jsdYtsibXt2ikLWak41c9y0t88n
ueJ7aoIulGRWqCne0b7wPCVeH65J87hFfel9122exA+n67ADn1kueQ/yqoXSOFCiBu2sIUnHIbJo
S/K7MzLP388vAVwRPIbOgVnw39ufu2tDvzdLB7SOsyPENtHWg/VSFBLhkIXzjQA/L77Rc9ZFPNk7
I+QEj9juxiPAW++ebLWxUH1jSTUA7ER1kAF0Al1rFG2irj+DdGytfbG7ZNStfHTKEG9gIVzdLMWz
uLhr/sX1YsiHA8zhYyUI7q5K5QYvmKAt6jj4YXr6HQF8yJuIKqFbieAjBwOtsmjIPR9dLUkF77by
PZvWk5w3zMzHi9WpaW491krFoGf0BRsaF5BqCRx3paMN8J5442Te29b46IaWIXE460K6DOCpIvHh
TvKz3NQ6O26iVQl0hXCWez9aYwcb6HSagWzPmbwN3oPmuJIF8Kq+e9AUk0NyCNbBXQznbd/lVPGF
+YYK1kngAtQiiYEBulrsOmpp7RrJE7eZkWFpfHd6uQCdGZKjS5jfFXisYxlzvw7eEfKOasIJxubq
VqecQtVsog8qsJ0TjfUoujnUnRwFhzv/vWbgeJytb1/ktqYUqdO6CRPBtpTYd2rKunM/4fCpG180
amGwm0/AXzGjx4ROVjO2mcOS4HjFKhLNedqbOBMNiqgJvek+oyS9Ij9OKz3I2V+TORXzWr/9gRGM
urya9keLe//512A+73fzh+9e7Uj2IfQxNnptR1XweOljP4eHGUVEMJJkmBmKmG1sS6r1oR0fp/o8
Cb1K07np2wAmBB+wJ0OM8jwfy9QidHoN3W8KLPVFl9iqy8ak+VfpjyUZ77LLEHseyebjMcB37plr
WQf1e/3DOnUBwf0uwWabPEb8WCfzxTaH9w8ReugpUhc0DKQerxU2Q9zLgz5arY8f5QQf/bilqhfz
NrvJ+bXCZCx/sDGWhTAQmF/4P8hU04zGEz9MnEgkkjmxmD2mep2pslr7uei3O4trG4l5LBu3EoJh
TOcSbQkcD354/OEHxYEAPdZKnd8NJWZhuAwQToAEQleMIuek+YLWebN6aLqlZwU12TNpxjiiyA2K
hbvLcUjJ6vLjQQLNoSUNE6fNR67R6w6/yARXaYK1sf9+olWzLs9Ap1NihmOeP9I9VVFG/58TlvfE
sXa5HBQeZokwzMvfD6rBUJ+dEf91JyfpkOm8FrR4jdwiCeH9VsSbRyH/giQX05FASZ1VsyLLINh3
wBza7fsyGteEcMwZTgsTUX06Mq6VdzfdNjCF0j57AOaJ8tb1MGV/XTFlCxGDVrNLZV7KZodHc3pO
3P9cCCvdb/jDGMc/zLhOZLvsN5QjJYoOc0j9pUzK3xdUJCKGfgb2FbVK05dbvvFUvGJWXTdukvR/
2+ATOtgJDLvC+YVR9ebvcu+v19U8ifpjHieC1KY5ZgAAhDormRSfZpu/uKwEgbXiQ0OEEHPkvVeq
z0zgyy4KNLbu456/kX+feLo4ZsVdjB3QUQhBsDfiMZpyHYsb+q4ZqFPN+HMIEHaE+YowSv58xzcK
t8m90upUGH7tCdCFctfY+g1smPMUOH0gar27ntuGy0Q27GpINAcYDclUrfhns2TkYano32G0mwOv
KuDjAz1jskI66ONAaQCJaIIynHsN7nVoLKN0/PNry2aLrQP8DCukv7+hAxm3HO00rwQCiVbqy4UD
qrCvkK+CmhpR92KUp0IgIWdc3+y4Lo/Dn1++baUazghOD81G/6XPveVMmSxSoGWv9DIbkr+MPqHj
VyPLfd/XvxJv9ZmV+BPuVrO4cGpiK+0bQnsCSydMNW3DB3uGUmTe2V0+5eDB+ydDoSFwIuPD+zwZ
RFaG49dxZAf1a6VibuAqFjsc4QOAnGhMffumsAujEobhKsa3HzHs3AG8Ku1zDnvniqQW7CvNuBLE
AuPJfv3UCCnk/S9gTXpIocDsBYFS0iyaKLLjlT8EAfXACMFwGzi0AkY0owt0WNSiYL8kcsjUmy0i
jFhqhsKUr0/zzsecQCaFo9ORyWgfnFCOMUcQjFhRZ2GnsxTQKRU6YegXyDJ11KVeKmvwnUQwW5+/
FVJrOiSk+Ze8li3mZopCdo7wpUezZAnE/3gu+8Hi68GJdJ2MpyGjBWBpC4QgyHdhB3l0rAougGNi
E2tWHlicO3cSbJv6YEu+F1R2o1hXl6Hre7PTYCM9hrOP8n5M/5WWQDDTB75mId3A7dixC0/rdVTm
rlhDj+131QGWk+1spSx8O+EqmEM25euD+PqlY/gd1E6KS3jUStIg2wN71Cj/1oAeSsJMCyXrZYz0
FWKxUSLVSzNkrnKa8iqsS15FyBzY1cl7TVhwNsSRFWA9iFuiKGfUh9Wmc06VIgdHrFa4P5fOyf+6
LueoxLfMJ5pxiVAZK2ywulTOFoSpi8/Mipe5oCbSWOFN6fAW74wh2f/YgYZx4YklJOXhf1TgQIQW
UBZr6X0AonCFSeAmCDAgpJytiZi1Em+t3hBBcdSM7bB6XgFISesaDYxh4NJnkhq8hMSeSXL4xNXD
PmhsBCAuqDjIstFVyqAnRbeLfV5HG8usxvCZNpflNKQwkl6HbXfNLupBpVNcXAv0RETqhO7mN7A+
ytZ463uC3FgfaU30VZiNc6dha28DTA0vKzQZUjJRSyaZ003JZ0AzlcdGKKGy+a5mDwjgid/Q9YVd
uSnWxOJ8jhXA4PUya9+iab8YiP4PNd32GjHY33Z7HeEogopH8zN4DNHQlxUVHKVfQ35HxsKij2Tm
XT4ZeOaMwcTxzZ7W1exhhGoQc+A++ozfaw0S4jAfkhmly/fj39btoEBniORwwGj+/EuhjJjOTfdS
Vzh1TewfxTIAd7/XHredE/+sIiTq21bX/SB49oYOQ0ghCdnPU8HYTSJ3rkDjy2vvana5bY6X9Rpr
FpHrObQZuSgIUGgaN5fIoHw5e7kKJNF0T6D33QZ1RdK5ta3glQK+9UJ2KqOAe/PQZb9ZK7Cs21r+
jNNUqGkap6v/XZOTqcNT8csqrVS6SbgoIhBgeY7A2kAtSoQ8fJtPd4kxAzwU7J/kFzdKvrckXKNw
5Y9u1d2NGQrbFU402go5FXR1L+IkIE3/LOWhKPevldMdOgcS4Wn6J0DyNqaiLTTbbLiufKqsZvyo
mPv9azi+Ig9HqoPsVQ1hF+TZUk6ewDqUgYhuVgRIdok74EcRqKzZ38uUXQikKzZ240KLh2Ij4sP1
+uq0nBW2hSUKbwww/As0icu/3nDFf0d2lYbGjk5nF7CIHaR4s3qQjvoVMKwiPB+NheDSGAJwp9HN
i9xioOYiLA8SYgx9duAk1Nv9wdm77n4Xe14fxsngXdInc03cFCDhRW9ZBxHeuXPiqFXPeDN0rpCL
PBqn9dI8wvzrInjoOluVNwcuKbNSm83tsdDoKyjZKl0XoSz4d1qfiivvkPdf9cm0Em/0SCNHLJvC
XSQJjFxkfcTo83Vk0J7tWbaZZiNfBHzz4oarDTro3PPF28eed8ykcwvN5mGF0EzhQ1mKpBoSWHKF
lrDQXI07GOVz+dHxjfp23ozLBTHhIUe2xKqtpaUeGPvTx22XmOaxJcsYyt5j/d2B9dPgnFh8FZtq
51CPwQ5EY8XOGnjoMh7wH0C0o8b2Jadt7yc/nKn1OP4aqGG4BWLAdPfMGuyWDJ6DBEOImdc3/cjV
ZMNobvJy45jLVtemtbOQ9YKbM1GGnVuXFDFJC9YsXHvbqseHm+Qch1b+d8qezSAlbHu/vCz2khl0
iZkxL/Qa4QeD2wsoGxF6B6rfbVBofF7BpFyN2WDWeTrAYdpfj+5UWsqn58AwMfSEIHjtor4rxFQR
rf0AvnkvtBcPnF4W/M2fvarMjahZoenvWmeNNH6uFqDl8LQG7j2/Y5cEVgpJ3BEN7Pnr/MFt2cjy
slx+t2knB70s9vD/5nQlkrrwRJ0pb8O10Eqauis2Zf5ZxhutEjo1Uoyd8vQZPKZYycgi+56zrgqC
XQbr4Xu921TcjYWvcxYD8QjttMYacwkxjZcdfJCawovoZaDuyqog8+AbRTrIjl0Pt0xj5zXLSu7o
mPtfMB1q9twIMlPktA5ugjrQq8un3wIOQue1HxnUuedLVQv/svKRH7K/rOxgSwJ81EwQItu1zpIf
kPjev9ggluTW+YWZatEzFB2Pw2MVcmT75DL9v1yL0iwY/A7Rfys6XFbPj9KPifGqaeHCDxVxjxfM
53k2v2iZql0Vc0gu3yuSB61U561fNcyxlMT/I/3HH5aLLb2OHmfbbXeH9yDZSW4jg/G7lH4jdcTf
ViBdq7x2Z6YuiKaz2g2nhJIn6VuVYgFUtK3gDYrTYFFP57g/rRdpD0yc1JjIPuD77B7JJmPolq7A
BotBlR4UO7mISwJ7VUxwGLhmiHjUkUvN5QT9DMcLBLMK9HSWTEd6TMYQ1gdbvDOU7TN7v5HkmzOs
eFOID4RFo9B9VF1AKxovGDpAdPWRAgFIAY35BlundhryE492MQ+GC9aUnN6GktZHK9S9zJ7qoSwh
cyPJltnIqC6DvXEj6od1h/ERpzlYa7M+xC4VYFiTtguUNLNJiXzHWuDmAYuAMEgPW8SSDropEX6A
rhnNe6X5/WGRfvVTJz/pdUURFxBbQuqNjlv4boQVWnxS3pAhYVupaAf3yuOa1dyDiKMlqzQ8VcKp
yboVScIRgODvrhfYzuoIqmclEIRNjLCMVndr/FO+4bRldTyJZy18Z7bSNmuVsXVh7EjI7oUrYyt8
0egZChgv7jppaAii52htrvoZyDRDBrNREP2h9XwpcE/Mir9QTaGoHu4B99xgaQ+216Fj+lnHdX0d
3iBgnykl1GXtRxQyBTmBBor4X637n20lw7J3F/iiMjVXyjZA8WQl70lPu/Gk0KcDEyVZvR6mVcrH
LAukpTvUho5yO1fP0eBiAu4P0EQS82K01svDhi87fVU0gIbwidKeqIxt1IKu0+omiix2h0c3I1Uu
3Uowcb0NGLaXVZPG0LsTM48+zeZ3JDM/d7KXUisZLYWY2yQWaSfwSyxpzBW0mut7jBlSeL3S+J2C
etPR8hgUUQUaCDnYaoLJPkec4loNk0gDzdP5ed3fHX7YUjx2CGorBgbv1oE1ktb835CYlPl89xYS
KYzpCud28DDWdtZckuIReMAQsgFEgA5y/N0SM7kVP8aoMxSx9z7+LUjuC5ZIDqWMLIfRM5qFFsoo
+vQW1x7+zQlGOrRgVf6YRiL4zJdylKkimmPePII9aNXzp7cjOpCbj5MNh57cFjnWBsly4wi4faMF
Ynti+KxAwMWbn3rH+z661Wy+glGp2hEqtkbGKWR6bOhicg19Uw75fpDCrRYOE1TmB2vTYb71VeYG
4kFkGhK7ad5W4nRS234Jq9ioU+k4/yM/G3BXNosdUfmg9cSPcKdqN35ap0s8QObYw3Lbg2xCk2e/
cADHUKiEfAyUYkDUj/LPTLAuBsnroA/95G3qEJK5Yod/0BFZFQSCHd/C73or92N2OO5dMoPO072y
noWMtAkm64jnZouIIBSSk4oygy9rZN4RRcaSr+VqHRoiNx1dxL6/a2DzpXnRz2DnzR9RNe/Pnk8G
w2YpBb22lCqjDDRP8W2+/afGkCEJuO5tVgexaKTHKRUQNcYmxCJ2ls/5X+A/9yVvBUQw9Fentsu3
btVI6mY7BkywtU8tNlht4jspIZ6ysa436ci2T9nwt0ck51YH08feuMkqCpFwfaiKIIXkN7S7AmLI
qPBar6WpRBbuZMOGBaXG27LCNepymRJFnE6yMgJ2jzQkTh4uvTtm8lTZ/hfZGKR/7IERb/3wWmIX
M65HLocA4G6Mh9ZjybHxU87e3cdLeMpsLur+3Tnpnjkikz5JD6612NccLeCUYX6dNMZBgz2GDS28
Aj3/bb84XO5SKnAJfdnePuBVw5GazDAx8kbNAu+j1MHox3HPBkbn2fbJKcVSoFTSycjpMYdtIh5K
qf/sgd48JfhATal9ZtPa+P9KudIGEM/yoweCx6l3at5elR/ZCpb2GNblVSjz/XWNJtUvnvO+G6nG
2DQH2MtaCCyNg6ugbXuu2oIagHxROnkkXzThqAycxKhKLalQ3mZn5jAIqcrjgKp2pFIeQSvyjqy9
OkWKZC600N2Qs50Ua0qqMSanuxUhVWiSxP+L+bm3KbaBTOzD/OvQ8Qu85kJYFEHfGmn9HqO5ZhMZ
RJ0K5qz7XZyTPJTemJnRuq0i2Z2rQuJYvzJR6aorzizR/2cQJy13uARSV5hD5f0/+uzRsup1yOJ6
qoC8XXhBJFACGwVl4GgpSPuB+Cw/yhhuvjwmjNO2yuERUxmsV8vXVXbXzsRc5zMh9vYjPygVbnYC
jZs2lzRYBtKsDAlaodjmN5O39jqcZqGwJNsXlKkJ1RAFcaO3/BxxLU82/gze2UqgorowE9+vUSc/
3j1zQaRmcIM54ZAusOSDsky97FygJH0ztsFqaRql516ykqFl+ALJz/BcpwOSDcSpzgRX/sRVCFl8
obr3jQZOoZkgzkUohg5nLRfzdfQ9uWSFIDA5l4wRS3MLp2ysIfIFzPzXrf2l/djl5zP+vlCV99M/
tTjUhSgFa+1QROVksZVO4t09lgnJj8U+Nzy3qwBRtsRh/1gUcsKVWk2VDIsRN6BibpNaImV0qGyt
P8b98VEPa2SfMqwf0gfhBdfYYozVy59uCf+hqXagB4L4SUupa+1rK9N2JHEqfA/1r3CqbYzljvnf
r3Vj2j32i9DibpqGxlLiRB/0aOvyy1HUQ3YpCNqXkEF1R9nd0BkXPl1UC2KGVp8eatccENacuJhZ
Ikib4qdxvHGxlW13dxWSRsUq9rRsAdbtnZnWjiend6QT9U8L1tVAL0nW7Tl6N9HqbKEXVHQWwRjB
l3U5LB552Yb0yt3dtWZ73309gpOszPGKnOqfkS3W0MiTzpgmZ4LCLZS9raEUTY+MV7AB9fVSitrd
UQGvL7PXD1jaODKNMr125e+tcFFOZNyN3d1IBxil7fLnYXshFTCLH0yHLF2tosisfGk8YrVL03s/
Ay+xu75YEZ2Vpv5h8VKz9vbtUPzSwVzUtRvP+fSvt72j3j/Z9CcsOrcbun0+9a4p+IKpKvm7q1WR
+SBuFwHPqB0zeTDrJteVyGeiRbz94HqHVN883rHr/Enamvu/vWFzQAcwO8VJ3AavPfMQGpYINgPA
2PS4QhiO2fcGrtjgPJts+PabbgnBZrdud0eEtJhIwb/Eay6Bhrsp02RyRauydk8hImRpY8wXZS1c
Q2dNvj+khsmbe7CQfCkEYivQ4uV5ny/zEXCcHzNGyWm1+eY2UzFgDNQSCDNUstXhc1NDvWm/ZQZq
QuGChTn3+wtBNT+TQOVmaJUtZXZNhMQzO/gq/7cRVJbuGBEBuPo/8mwG5LOva8+UVJh+Hnhvrxwn
VqoC6+ZEvuttFJS46etXCFQl3QRwomJcpCyUtjwFTsjT4ADuHwclMRayATtW8N2HeW68pjE6iU25
RYe6U8+dYOV/KMH3sbB86iHJOy8leE5t7qXERlueMpprR4rsBWEbcLTNEtaLDcPCyPUr4WI1E9D+
rToRk6s1iO2vg7xtYBpAc3uXupoeEJhR7JMMjGGtCKStOSPJzwkmzpqAD6RHkXg3gNtF7Zq8/Btd
Fm1PiDosa69IlA64sRTb68i86rbBfDjRIz3oAUSmxG1LJ+CgV+TcMYjVAARgk94eVYwd7ai8DT2h
V+fIzpwXRMMlEGlSXUJCw56yeaXOI1jmM3PgmmrCf0mDFYKDlH64rGXFNLXfXAxbCspCExifXMlJ
scv4mlzx0ZjHSNyAeclis6gFbvK/1qQUtMMd/IhhtNY4l8iq83tKgCxfw3zL+jDcFAgMB2HeXvQi
szyh6SPYUSazTXohNB1RFW2/RG4dhplKS1i9Obk/3sBuji2TBW/cQLdczpUifYod3f4+5JysCHwy
7+5p1hbBU4GqB58xUnHxTMzp8H3QO3/id9L2IonjLi85w88NsQWYGfZSQApTmkTDTGLancSS/cgw
qYuQoqM0/c264rga7+u1pBxwHU3swuk7yyoShox2/DCly27plTokBrZBkSIguFaCTPemPu+5Cz6S
f5Hx52Mu9z3dKvDtQl+SqDW/ED3rW57iMAckNx97xvQIkiVOkJXrF4hOoGAAire1p0Q8ovwcMvUN
+FKedkb4FQBKNy/X/tAVfvvNCOTK5aFALLlXsIzUIBdqegIrKnFu+u1vzZADKoiALwWdVqxhk77v
OdsFDeDd6P3kI6yMsUCYd0nnnBieZfTvZFS6DRoliEAxiFCocHSyJhghnglZexcUtRG7AV/vDUlM
teLPzcthOHvY7m7l03FjfPVDMaXAwq3A1Qla4KEUsOw/osiGQuOES6RBby3pawQnAbFhy0D7PgNY
5NFY6z195GR1nrIJ9QJ2HPUFh5f2l3SGUbxIYgLMVPv1pfw9KLGp80lBmywXUzKJ5no0HVfyHAzv
p9k2yZM8gVFBsDU9pOrrS7hk4ELP2OFJdi3JvfHY9DtSW5XpbKoBcvj8UrPPtZekzfN9RicS2crX
ObX+uTpBZPmGfeMWoJIaniZs8zhL4n8sSWeJaYvPLlOOJVDPTFeQM8iwxrB/Z+dhOxEZxIJ72Jry
DxhEHLwWvtoGnuM2XnevV9SkY2dQQEnTtaY66fwNqvhDQHW6zqulsdH4JuVvXYRe1plzm9nxYpbG
Sm+BW1r/3hn+Tq4VrYHyicnsOM5SnwThPO9+/18Vhoz6PDm5zjk+IhrITTD1up5mrlX7X7w2Gvqs
1JDxSy3xTCES2YzHPQs+UbtU+5k/lPl3at9dnpyw0wP+sMC2hV1lp0PK7F32TWetFQmCMZK9iGYr
S17ux8PZH970YRfuWwPsTQMrmXtZqONBQ85YnAP2wxqhFdGfuOg5aVSg5GSvhs/0z7gqiTVuVbrh
qjNfCB5P2q+GveYB/ksbZUVkq3PHKL+1JYNJJlR5IPi/OYkR+wPFbgEt7ZN0XbQZ65LwPqoDdb9Y
T17586uTqODr8JufXvgCPQEgI6wrkQlOCALoQmpbqpyz4XM4gWeDGmAiP9rBOqqPQBAV1LQ0vmev
cv+gwnr1Sj1q9QU0+HPKa/RqaTUpdWQIcRwkKWXn8GS++eOvjUdc1+LkilZ86sn3A/yWhQVWJJaD
uxEt/gVazebOVAdop1Y+hrktWejwrOEVSGE0HlK23KxdE5oK95JwgF6ahYCIJMiFac/3ZaVdj1/k
pWW2EjduqH48Vc8GGnqg4ovi+QhaiPHrY9KrZ+3f/8nkvSfdXBRo+TR1N95OqZqBnHzXr1T2uX+t
LSXWhkc3znySqBEs8OQFuG4m1XSQN1y8VNUScKwbIky2cZ5p9ShYKbdJwEnS6gQJcL4AwkX68jaZ
3C7gv6bsdrxjUbmybI0UgifWK0scV6Jy7HijEpgWFj+++C13RNxXvDVIkBjb3byypl8YbmqUdsgZ
+Baxo762zs7H/J4T6hmrJyiB5ajLjwwceVmXu1J88ALzOEDZZ4GDzwaAW4f3oMMYP3nmZTGewET7
0VtR32wJQTmoGT9zflq3yfxoq97X5vsKs7TAilwoyMuueXhXNz4GkBSFDzo4I9fnAkfR6jwHXLKr
XRJYtlNQLeYcbQl9c4VJFvt/4Xo1tLyRuPBiFeQPd8VuYVtNkZvCHclsRj6Z+I1Ign7ec8ZvSRX6
HQNFFeTU6V83F3JVRjVEkCZpWQCOaRXqpZIf6O6dGo9M2dQ4eHVcDqnAUhb4/guACWi4vTVV8LBb
YnU7xnPoIH5bRd5nLBKY9lJMapBNrLB8+QsfV5INyXn/N8loj3QEtXU6D4ny/I4sZJBjJDxjf5KE
2BARsFLEoZ+xfxLOVckjDElEtUJsTitBpRyFTmcyZ5GCgq1rcw2L7gwl+BF584a5r7eCrBWH9Hll
2ldIh5R6kmkqY9XvAPIE1hVzkKZkrYlqch9ejZRo/xZtxPYFARDyC2HRF1ou4LMPsiePbtw1DloK
Qmyx6j1Qxrz/5pK3yqoy3GXltGL8QvWleW5By2H6XRTEwePypkv4hxLbDmmP/ZdQuKYozEZQoMsO
tyNY1YAOMr96ahNpNwsjlQtcFA7AuDrr2VsjbF3d++7vcdZ2n7MK1emKMP0qMS30U4pvddfDVSoS
tcTbWdiM54PJ57kSDl2QYS8Wv60XlHaQhm5tDWQN2MI8L0kRsLlxU4lyeeV31sZta194vkD5AzD5
awe/Cch19Yb8+F1UuNLBD8Ct/Uho9tSE7Rw24fURghI4JgQHVwCxUz7M+KsUhez4vezGnlvuvmqc
CVyaOXE2pX99eSnpYryvYn6TDekRh7/4vgy2BJsSSqtp0od5ke7tmWBCo9TelmENZJmE2YY83sje
e1tmZOFoMvCRl2t0iIT7Qs6/yO+QAik11/4p/8oQrxGPJHndTYALtxt2FMx8gz4k6Y9MhbWF8/x8
TA4ufGUv6HiJURBeZHf4pcs/yVIb6ZPyiW5BDi9xpqMgj56g136XYGU5DsG0l3qJsrafDDAUjx0X
pSBDBoY7VslvyQUxASUMy5qiSIbtXpm5nlQo09emjJmDzRtvkMd5NCEcG8ceF80FtaLnJxBKNhdK
pzBnzVPXCQjIRz3tIWHaLnDtABVC7e5O9W2u27KOMOq5WcrWtyKjyZU9ucezCu6bD3nVylS5fnxm
M6KWwBYdUXkoYK5op9TSbHSsxkWG7E8CrKcvOjLqGJN+MIjf9bxZFfwJGdjOQAosrkjVlpBgPxds
2x8OGiehVX47nx+zZ+Rqqz2SHDFth9KJqPZ6zyXf8cYxlvuh4ghETdF9O3GdfHVnfodf+AXH5Ril
Me6A9pS0FePn9m6rDmJrz2xPBFuN67B9JnNN2WuwCcl8zSJ73JL3dZhjFi73Jq8pWhwBoAQo3kve
tTtT6BHBVB12Ai15IxMIRdPZEd404qaEL3yHXZY6mJzuCqXVpE9bJntgMBe/+oE1SSrC6hXDzT7l
LjZIDgEWWVtxrMQ6HE+fLp43/1r9bEVSoNF+a0DyFeXiHNhy0mCN7yp8fPG1fY0z42I9jLfwYh6z
YSQRbA/Od3ZL9LXezJEWzPCu41kNN+FNFV11j9eXT/qq5V4kbOek3rwZU7I35gbYA89NotV6jV/y
7HrtVQ9YhIccPzuzOcD8XIQyXrBPP+yeVE++D5v4TZezDgZ1Gtl/YkBbreAqhHjMr0cDmit8a5zZ
UldHt5aroz0mMeEsqWeiSC7/m6VxOyhN8H2IZtoSVyQC81SiwlIDPpuZ2DYqWODDskYNvCTUhNMa
cU00Kq/P4cDxy/a+QZnL8vkSNBW/5MkivVZPshaxZ4qjtd0hY+nlWm2dSUgxjz4c/dyqn+MKmE6M
jD5euNxLvWSfeVbWb3DuvMCRQ3kJSCVrcIKQ4ZLPj+GPasxNubMNbSy3yMcCe+QwVO4SgYa+S290
Rws0moZY/Gni5MD5zjdqCH44W5vzf+iGhu0JtaDBPZW4aZ/C4qZIUUZX0ol1enw350Cisc86ZHbC
yGfx95yDZKDbJj/+nbeeOw/i3ziUDHJhzOQ0QUW1AotcKfyQ2vglstB3DiRZ7mzzrJ9lTfo6cxXU
IhXlZWvWhZaw/aHAOMZS5PzNf/EbN4GRbc6Si57m/wCEd1XeKUGpe2zOBM3PKG9bc/zOzg+BbQWS
fdTteNLb/xYWvGPFLE2GjQeekzDmk8tHIDc+YTXSozOuAFRq/c2SAu9VkORzyWCDSnEj0nZQ+kzz
pqSpjcj6LV8Ih+YyD6/IJYyw08HRlhByFd37DyhktC/e0wS9nSFoj0wg9jCglPsNTe0gBNHgLN2C
RUijzjjdwFC+Pfxd7cqR0OcqaG5YZoHWHUJIrOqflvrA/OTP+stgodDkz1UaXST1XSKNtmfRgTnZ
SSP/3/SqEAGiL6E7L4RoOFVzepQJvp/5PSAcQK/WeTOVTWKvKDJ9R40tar/UPQ9UeCbrn47vEG0t
WvKDD1ccRh8Q1jaIF93chSv3jsdYdd+ArGko7vxSooUCz8AHR87OGzy6FALANUBM3rJDq8JAeyJc
ZOfCnLMQ/OJR0Myr+bbJLAVY8jgRR94IsxfWBpV8URDF+0RwQu9buhm/q8ja0rmpMNtSrS5+CeKl
+FfBZtlrxMZTbquzCOugQIXsb971p9w1DglSGrKO3bcWwK9xnVlhg8KTOB1lLFcX2ZdZeq+SKEeR
3UL6ESAPskA9G7YyqFS73ve9KwJBr5dV40hpHHTCxh1XcVlQQYbxyYtuO2vQbxFblpk/9G2x0ve4
mmh5mqK0DmXSwFoJ3iQajKJqp7YHRdwTf0Xzk3efpYLjpFzNHx4NbOns3ZdKJhgO/T/Scl+1MWrs
S11QQSZ39d01UtN6K3oED7zG4Q84E+sjZI6XnqSDfiOdj5HPHhIdEx83iSPUafsx+2iceosJootm
euMoYz0d3qx0L8caxWg8KrhwknGZBdvKW+1aC9Z+xRhFDVqL6Tbw0G//QZGH1Om+Sg3p4a1meJFC
5YmiIFj/ikij1onIeRXX3kYGalqYQcy9u/jZSEyFFl57tQ2CMfTQG5VSeF8hhTlc2L6Brn7bAfMd
O+ZSG4rZPr++Wa62o6BJcZGkMqnxLz/skHIkhgKO2CuLPqh95BQ49bxHnDe8ENLrcfvk5H3iWkeR
gmq2hw+d+yF51Yo+aSpCci8vW9SJVBevRHd6+lcSZshihpHZQfnjfatigpjIVfVoYYWdC+ngxg+I
mrP0Fih6Vz1WetR22Wv/P6TCky6KBNIRFdibPJ1D9Grm2JGw/7RXR1557ZdBfpXvnLBShB0wIlFv
0P7sbeVpNP8uq48rIU5LwKA4Z5XA63MWGc+HL6ijJqrWWIj2V9Xdc+ls9Bxbxss1BnEkfliXGQMK
mTUhADFZNMNjWimirAyfrBSyiPN2m9KqAa06uBcu66cOjuNQVd6U4OC5qhuxjAEG3L8vZFx9tbDY
UOnEgOO3XdrQg8bfSWn3oV0TeV/MbD99CcFcQpKAPrdhF2e1YCIFYYbZaqtq5VScGlJmupft23mV
PlJocpliOPPrMLeRLHZvxHVzRTb6vBN/6X2oqakMUFXN6ZZqhJhqJyDhlVdYexWQuTz970rTSlu7
FzCP3Ath4lgzLQSwgpgD2RVxT/pKETOnWXXPNXsVBWxkp+3gaCl8/oAWBmmdMQ9yzbF2WO9QCmOH
q3r7cClPMgsiHI+hBazoua6Ig792zNA1RuDPQf6lkQdZgpWOsRNC3J9tp19jsa8WtOZLkiHL7vAH
7jelzIP+ToptfX2aSMiNWIq4hyQIfH01ZI7aSaudWcdgJryfhynVGdY3TaFShfmdghOZ54CY4lGD
pep4PmJgS4QjQuPtxAjDzH3BVo8692rWvwrKQ5XJOJLOc1kPZb1MLFu7wZVLz3wcgbT5eGL5+kGy
SYlWlHVBHe+dZxX/yjvJ37gijxLOBPpnL9iR9/FwkoKdjyapOd/WLB4svPW5nfi/uVSzrwp7ElLQ
o7ieYvtj6q4CdLVGUHRTGqt9AfC6bQzZWnbQK3ibOMRL1h0rLRd9kQu8wbPn6tGnQQ2rkdW1c46m
5DvKHad+jQ45TmUyWPhP9NRY+Bje66amL/0+eOlanVxQzoyfP5Ivp6zFW/PiqBtGSoPqgRmSp8eN
QJCbUkltaoYyhpXhvTIivNyDtbvUc4dfvqP2n+XAJzVmEZNWztnXs/v2Vo+GNysN6Rp+JTHqYrIH
hqU6Jz5igBM/QUdQyn2wrG2A0MAe9gbjFbRQ9LqSNfBR28fdhLJHpFOQHa4XYNmsAgGlLwskgEcp
oHqJ3JMwtgFXEY+TXuvmyO1P+BUvAKLfLudZI35s0c0yPnsCypEkg3/B2uM3pRoUtrweOTmTOO/R
Fh+cvuUBrGZvwI3g4oukc/sGUhOjOdyTjbfSt9Hh6tFZIQlKFg80ZKxFmeXcYptFV3AvGZeXGbQK
fCrBn06Q4HI7x+1fkcNot6IhHutETZdkqP+WE3JjAJ1TviMZ4vvrXHFEQDJSXqCCk2++QQ7gCzgK
UOdh7R3A0o5aw47lJMq2QPKgbLUQFKnqXY5A5pAF11jl3mU3p/wEhIUYTsZ7oD86qRINnseWYBuy
wPWpZw9BEY47sgw+bS1ijL22oPPpZLqafUDZf5jcIefCE130NZprWbIQ4hI/1GqqoJf0MQMZ/tSV
+kBgYeysOEd+C4DtBxFBVqMuT2YMqXk6qzNeqRdF7389+ynqN4/J6X0dd0wXyls1WgdKo/4XOJuA
otVsDKhH0ACo5IYyHRpQHKOug2/bnzyyqvhzq3sQdeRzgpjyP4fkAZ9dj9E/0oXZgAclgz3uGDnH
dvW5SwK2CpdwecsW/LAZ39Yi3VtsboDGJhu58JPHzFsUcvIw9ghQk5u7w2xr9+f7zw+yP6j3ytIj
od/p1p0ThZKa1eyj5sowGN5NCpynYRjFCTJnrmldj4p6SrW+ff9DkBt6zFjpmUafrTUiioAGGbnn
Q1HqfrVlCDl/fZ3P0h/BKSKbNNt3RJ2DjUcXpwTk8Q0DOrb8nRVfi6KXDigH1DbYuSY/hGRMThfI
q/qhprTEoNekMN9gBKAk5bmg6ZV8i9MDSnc1OrrioS3ukSBtEM1YnEb3pD0iZYF9m/Z+oIYM0VYC
P+LFvFdQ/nBRBQh3wMN6L/F5k7k9y6/i7NbNeHF1dn0goUcoeGO9M8vockPXfjJNrNiaw4TVoH/n
d43ctsrsrKfGVddNHeKr+/5RKuKroGntYZHC+XwX1UhO2ZlMyomykVFGdyrByXnsyFDx05u1zDN1
88Wx2bIdbdhljwbqPqh/pmuPl65xTeAHFp4AC8f1joSOMNgMejJR1obZ/hb9HGRv5DZK/EppwR6B
ADDlDa2os5V9eYN3FF9ymkN87bYd7Lgp/YpOoXDU8i1uk5Si9Vd+YS8KgCLFmoLYHXup5ve1UDpk
7qdyIUu8NXAslnZghO0GPi+Xq9qBAsKjKX0x2phiFwgQZZf+zr61ueCj4OXmSoE195deQ+sFbCRF
QO+90mpj55/23jfO3QwIGwoTqmLB5xvK26uevjskfntxyZHZrLuFQmhuwwwUHpnFZfw3yO3VRL4b
ubGF7paU7mNkGnWkUE6bQt+XgrvO76rPGN3MJ+vw4YFv7dKB7JUQHGHx+PPxqbFAFIIpFLZQX44o
tydQM0tY4MjOqYgnZcQ8wFtQea0EUHI+PGFYVUF/CNmHDkyUw4KkI6v5o4bhQzTWbAh++eeCv1tw
I5mhY/J3UwzO0uCpYsmH14IJclt+X7iAhJf+25svFMv/rxPfA6pk0y42DTCXM43W8g7YJXvXzVRc
BykdK/w5gfhTkSfK8hpQzAkn/zTWZk/di18hcNi8DqGA5puNlktYK1xdDGcJPCypHxnj5W2mLI5l
EBWQGWaaoUbaEEZSGRTF2lnjxv9TfwYCnbmEA5XS3kegcpzbsqVe8m1WhGXBWzDYnStR8bKhOzRo
cW3+/XzxzbBt/T/3IVJKbsnc2qRO62pF3RGTSnRLPESQWrAn8yKFeToJAm2vuoR4pgSi91LZXKeA
PV+VDBKw1y2e5tPm0lPQfgG5/zAnKoxDkIkSk953PBqBEq4E1VxYurFZcp2LBk/KmS4CJhp8QjBl
hXWirX9U9MilCRzmrgt9kuBT3RrAhkl70eBpQ4QufwOTRymA4bJgRF1ByDo1B54ZBqYj+5UtuBcj
p6bOzTB8bqsG8/BD552jbZuU79OhwhczHzKWj4bI5VBjk+MIXTPo22JnRU913qUTwPuIOEwOnQXN
699UxtgDRHNdTXyRDY1OLKOtzuL22+9/0G4ADwGJ/0sPjNhdOCEjl7IPrJ/LtJqSAxEl3u+0fVpt
x7EpWU1yYnvvnHjC1ErtdFdtutkzISBimLk96zHv7Bj8fcrpxonCB1Sk6Jk+HuNinJYzL4qseFkb
7bMeKD1uhJAyTLCt26z5101XfWo8BSPLYXCWLBRfpdddaaHeJdG0PJOlS/Xl/voGqYcs0yj1B4Fw
yVwjIbxh2WjZ2FihyDDITUlvhL9AtWU6qafjrloEstAiT53/XKb8WWhNj650d3FQoWcQLl4U2ZJ+
yWBVG60Yq86TZfxDd9gkCqaBmraC3lctowkYvUuruyBusHjMoqckdT8xFFoE3t6eJ4GWECSS6gEj
GKpbWrxmsGSUyvB8YIGntl+965yqhhk8zHfZGLte0x46FFU5bx/l+JZ6kT+MV4WDPOTeMzMyJSDn
aSMWse+syE3xjb1Ri9PKtr/rxIbBWHoO6YEDyxe3jBG4AJhlvRWjx7kFRrBA4YT3D9u7WKGerys6
O1w84N4qLcT0RSmZrASNBAe/UcAwDyGbU9twvr9/7HaaZvA7R1Tlh8DpUtAaVL4/k4uj6awWwXUy
H5Kk9fq2a78M0qwgkG/8ie3CwjuS0x0MFwVcVYPSGosVkhDRHAHKJkQ3FEDv1SJ+/lsZowWhJ7vh
PLn12gxSH2o3HNQZSN2n62wWcqB0tAap5B5PLnS8js1ZmX/sreyINeBT+4CnK6W2btFlLvves+8L
fEO6i9xECorB2MRBed/jzcTgTnBxXGMAvgj0itiml4x60G+/g2QVSpC/7JYP9khxQS8mZrSDRG7c
HRBNuWjVgluidfRxkWO7uO3oeUG/4XxkbYgOE1GxarV5fbhwBQWzdVNOSwPcXG2ONws2vpTTAHH/
r/68qx02/ySHimCmJQlnbsEyKyPanA8gJTclfazCp9/lEA1bMRCWS+jGf7NHuL3A9MQu9WpsUsxQ
tLALlgMQsyAsRDrZWf5sKvrrrNUptddkBnReiBMXgLZIGW2zcUcJD97nYg58wamu0AgEU6r4MnSZ
iwv72FTpzsmJL+6MXuRz2gGB2B/l0VMJxVJJmsLp0Y5OmU6eY8Dj3OQnVRS9/klRuytVDKkeDRLK
S+FeqxnRdM/NJUXfP2FAeF2Hl7gxs+qQmEhanWbocMWMHPNC6N3buFzxdUvNkpFWkyjrr3ejtF5k
TEKzO8o85yeKIwOTi8mz4m3aIXD5NX0GoJsG1EI8RlodFoRgyKlqm/mbjPbD6U67tMcMcgCTQN65
Z9ruAPM4xDNwIyda6CcrN4mONA2JdRu24/VJqp5kSonUMAHF4tdYnuMnTzfeBrvFzQgE0786kQH7
DOtR+hEhnvk+F/KJ9zZQDDGfsCP7PYvSaoHSo0TtqpZPgkJ/gCtM5nug0w7/ZS7vjcAGqjdVCogv
10Ol4eb2VEu0Nl/hCohaJBa7Rj5Y9o5tRgdWUwIeIEq0X3ajr7YyrJAesKDOI4AWD3gMCjeiEwV7
pArXE3QMxANBldfA8AFsnf8hsJ5qjUFaA1cXHYb/7wWa8is8Zms1I/5JBxRGNLxk0WUpXFw4e5xw
eGctqy746UTgVQHe60Rew4i02A3zwEu3It/Z0ZJSg+ngdRaJaIM73IDmZu5UydfL+xsvqAQ4Wt9m
5818BWkK3BK+dFiKZm/zEuY8UATIN3VwLwnohqfTSTIikCFVnQELZAiAFDN2xaZC1tkTAVBe1o+2
H1bY5CU8phheUa6sBFyViuGQpXkvv6uEpHyR3TWoFTbF82mP9l9/t4zQmGykIMA43YTND12zWgBy
iOUV6y1I0ddspwVhKdbDikdVoDbJA1I3FMtgHmJm+wauP28jYBx8Vjnf7Zk+OJLAH+kqOUQOn24+
YAPF+ukUwTBfW13bfNZhcz9XmIu2/CxrayE7S/aRgYx8kP3ni+GIxsirH9L4ixyYVfR/3RYkl4ir
ipFzky1Q+/s0sHsXzhje8ZLt4TMlUwAbfYvIa7K0aag06gGCFgN+QqwtmxIugMKCfDc/KegjyAQp
DD5J9ba0ZpBHR2qznt/High0FH+svMYPS+5OPgjGuUzuo/nv+9XEwt9KkeyOeCwIy7M1ktzF93+e
Cte2iV5B+Ncr9HPgVthv0u+FEXWgZ+pZiG6y+MOp90RlIdHl31si4aeBMjrCVTf7vzKmeIbfGgfe
cQd6RB2O4yhkij2JYCa01IZqLPOLjgw3Xw0HCF9i4pctu7QbJE/FQ3L+jRPjPwPuQ1GB6oHyNId0
s209EznTTnte/7hA/x4jSjTlXYxNLxYTMMKCammki4Bl7QuDzm8W4HOy7V5GR6HBWJ/8ieU4KPa1
Zp0J6lyJ3GgxqubZRFV/kMci9ZEItlLSSeESO3YsWe4Ke7JnB8AVcEoHfcXVfFOJCcX/IyWHDAmv
PFxq6oYJ/7SDPbB+PfEas7PBO7X61q9wewxwwxJcOHrKJJyybrP/JhRKx7XF7ge/KXHnd2quPmYZ
p4HAJa4M7gOpBE8tv9+IbzJxylSYaRxalYvTiO+8XL1T74SgXPw/R+W5Zm7tGySzKsY4LOWNu/eR
RRjEunN6QDk743/hvuodebXLVdsVn8R/7VEwV6IKlv0AXpMso6ppS/aKz+c+Xs+GFztp9EZ6iOMU
Jj2xKzUeKu8vfb2WgAKI1Y/Ewa+9zBbbLg1yIOgL4qAC/EZVJr4l/sqn1+HyvWBAspTnn6rJOjZB
qAAvaZK8G9ME5/mQghehlIfFCdc6/X26N0LdyFNvNlKKZJlhUC5zuz2LBqMLNagN//uYL3FkbED5
NK5Ul3SrHrlFQET0hOMUAskcCMZ4nA0mEhcngWd31fNYW8GFTjMEDsQ1vOWQFHVk+1M2ZYf1Vwr0
zpEshxtzoU/IN50A1y1bcTRY+pCsf5UAs3WsZXrsjtSPhlP0A/GO4by4eUyFRKpBrBd7U+X0fUUd
XwuSTy6KWxceRVVnDo8nCHBS0TCWYjaCJf2rbebMwIrSrbsvla5SC0ypqaBelNTvIuP6Sk0jUfHN
Ndo73c8lL2uSUFilZ4GVb79IG+6XkA5TeP468M0o3s46fsc3LKXwbqR0iD5rHTZ93qKC4JE9/+OT
vH1Sz1FlzCG/9Ebdp3SIGYNKG3bjCoYIe2APIiUU3uCRxvwxWJfErkZnd6BvqpfbnGCT5h2d3fPH
jQOL/lJ3OktTBToP4v/14J9u1iR3Hxxg/0UD3xEuz8cfPGTs/A72Sohuie8yxJV8HAnY9qiRfHyX
jQVLlIdUmQy5IqeJYDoD1PQpKvuYG0C3mNjYX+wWqFbdeROQGLbOHUxxzqwN1U0aoPBMAXl8YLsE
4Qo56C4zChgPJT2I136ofyjxKEF9spRRbnTKnNkamyVHkRXbtSt5hjOT03ekxbw6BFV8fHgdWcWW
5mz7TBqLvRbdykMrkJSntT1gQjHZQVC4MQ2a0yowfE9k/r+OPf9VEQfpyZMOIqQaAE76pMRJyIga
3eYJuwMvmPeXOv1Mdg/EhZo9B+bhyRQimc4ZrD1EKPTKpxOymfoPfOfJoVOXJ7k2dmz6ur9q3Q0t
ZZiQ3qVYN5cTCTHtRwebXiVS8VfpIlA/+nkvWFxXJgz1YWNZoWERGeWMlTKnCsDv43T9faMbpodJ
R99Xdj3MJ5NBSGFfFvmEE2uCVj5ELirZkSwOYCqwLlZYefJq/vlruK3xlzhLxL78PQQp6Pd84fcK
7PqJ1V7oDj54iqm1uz0JQTmaTEmMVhzVsGKdO7oI6izikc/sOi8NJgaLEf1KK21/oqEyrhQ+q5Yd
Wtuo9+8yp2XmuZKdZCLdPKi7PKsWbD8fLgOmKq8zzTi1BMnK9ZAXvaSoZEnT42tu4Wu4vv0mzpes
B4ixojhYuoYqRD5qVen6didcs3kHuTLDH9v+p3yB25+l904HvKOEPpxFjqOqIkg1P//Q5L/Y/pGn
F2eJ0WO49GUx+EkmT350uLYsaPDM+f3I5/EcNb/n5UynyN+EeDYxORcz2mJVK/8unFdC++SsMYZA
lvWO/DMZJK57gnUll54sTUblUDLtkYCXaiDzbxf2Wli+O78qHQKVOXbMPJ0ldhlsele3QXsrxh4m
hTrPbuG8Xnn1zjUaA7uxUF1OHuHsDPthg8WsWQw5bBDWt+ljItiEY/2s31O+7XIfXstYCRSUDCHQ
LJnalnow4mQN+PVmhK5Pr2cfXn0ixflIvUtDvr3oolyffdOR7XtLVY8oaMjHBfNxwnW0jqBm3Fij
4V8mdCGftwXD1/WjBijPulbbabY9oVBolEP14m82w4rFPPois91OISJjRgh0wJ0RyGwF0MXeWgF9
+9jmlDHSRH8qI8vS9yBZ5/tl4dFGxzKJ9FNlwCjyP8ZUy9gBBahbwNjwqn42vCfxGsQY72Nm0sOX
sdiRhZlsGUekQbpeCzYcA3nYvXiqdMpTzu3X6rBWhBcWxs/Uzo+bbKxt5XnewGqoQ5hPNiEgLGhp
2jbXeZ5EjA0fZfVrJEi/1PMxby54CgGW3Ieuxx/WN3qZHXA1YTXeso+tcE2VRlPfePOQ9s6NvQhM
6dQSKVgLfd1/yUVzbPE1EvWdZ0DTzISKsES/ruX06rcAW5+4OB2kWLjUoUOJmSEzKOwP3o2UjlTr
QhGa7ZX2nMPRafTts87IVBXE5sDAO+b2eNR2bKc7h9LQ6KItu82Lj4UZj3GEW2OWu1Jf9cKyPJVz
NlPbgX9J35uJjIY/Zz0XQU8Jfro5j3UPrWt8lGsyIShhUZNmREvHIwUdt4pybd3dw1Mz4eZu/AFl
wrjSZUq40M5pE83Rff+AjsfuPM/IEpyvyBqm6GtyDHKqU4CpTN6dbHussH8lWyYwZiXR/4h6z1Sy
GBzI6fPV+fDtgblV8hbqtyD8ccD0kegaz1mIOm09uaNEXtdT8hV7PWb8yFneMqGZPtGdC34AxSVJ
FBNWzKF8MSI7aop7Lrxh5vjSRFDE1bxpez6eV5OBcxUHjoG55gtLp0X9mspPCrPt8GhbGi9EuJqm
36dqhjdx2nOgzmd+o9VevNV/zyFaxcn0J0czZDy5tabbLfPfd1iyaui9mj9lD4aGSUD8xV+BFy1Q
XSMPBfvfbd3Dlj0+nrJnUUJGq+jBBy3A6kBT29HTjp3upxRdHwwUoR1FNFsYikd72olLITVtCxk/
WqIyrSNbR23M6wOI3mPoo5pGmRSpp4oFhZ1C0PPaJBmw8FZwCb5eRV1PTZB/qWIOAteeLKzWUw9/
Wsu9h6QYft4JKlmbICi/Im7+gf2LxhYcv4yobYF5LZfYFbU20WP5nU6Wp+zq2GGmwtZQf/G4OIdA
SnrAeDtZ16u5YJAV0qnub3VT0CsgFrjmdvlwsFGW1IWh4YZZAXS/aoMYMExMsfABmUmlLEw5l/oN
pQYyK71s7fByQHdW0lmQpF2w1tznxots2TWjCsG3x44biPfaJMLA5w+aQU+50WPhEefYGnKZSn7z
JaPzxv7fS21tWUtjID8tSBX8LPSPiRTaKTETu1wURBvQgPxRU/BVz6i/7f0DSCegtjUHFg7Z+g1y
Om7xmyBaLluh3aBS2q5t3phvasI6H7gAnNqEZwXjQYbFIGPDA1D3vyk2CGn/C5GQFebbSwQts1Js
DkCmLcF3VGm2nlPUziBVZvrCfvKspsR8Z2/ZODiMJCUiE5gAlg6Qnxsieu6E4vGhz6KpjJGcSxbi
A8wv6Fhno8Cn9uDWmErrOgEAzqv+YEp/ZkwKA0PSgzcG+Y+uHPmNBzLteK/6bGbOspPeRpwh0pHJ
OqVyAiylb9llCkgXQ8Tn4puCgkbqtL2SzCuhaRmBzlC9BT/3NvI2/1/gMT7VtOAzxp8mlbfxxF4v
MD3s8XBd/XAi1ITOg1EfCVV33145Eoxvh8eiYpd41IWuSsi8qKvU6DRKkCqV0o+FzL6ihc6KcDQT
kftg13I8oEOt8nJtb3bXoKfn+ouhXtzFzkwLmndsJigqk0/dxLfm5KatvK/qLJCNGV/NYwsHo7hB
HiHa4grIROSusBDsx/79tfa7eiAFFmaUQ94vIaaYGqsWubURJKYfDblqZXQ8/4Jmx+1NeRDwyt2T
L5ed0XrazAInE/daO4SsyislFTKtTTT8sevjaS+JNRyyM251HtGkkV9iMxvAWs2S3ZcEDnyzIBvn
+ge5ukaeyzogPLT3ehgZUwkWYuuj35LgjiUze9gScpe8lrCAKTEqaJFb7MI8OI9A3m7hBknLKcvI
yexEM5GxGxX3kuZy72547i+to96nqOj2xOHDzsBTbDtm0GuRLSFl3vuisApE7wP5m6KO0p4Y438Z
SRpX+wpgdZGnVdmJU4PZkuJWT4pnJhy+T8Gi1UeD3mxXpsRkM4mxf4LsdSiC89qfjvs8O5GclPe4
teING17BgFuthH1dduL2T+pY4ivhRMK+HgOCJL2p8kBSU6gBeTaHhQs5YwxHutL71J6N/uaZhw0Y
17nriqeMs6HudxpMMVrxtXJp61LHYEr7cJY6MDwfGqatLt7QDSXqISN2dRlbqHJlvPAqjdt/8RKO
6KaajE/LAyl83Ve6j78P0rwg9cBx2UX96D9q2cB8UBcryhlErNQqhVagIUwvvjtLkj5ZPteeNw8c
RLca4gIkQ2hMlueaNpgjtnICXYpS1WhpSxNpCFqChVWHkP2FL2f8t0B7GStmwNz7m0M8a8MygLj6
Ki79NKxwnku5W0qBsqe9Bl1j9rffvLKkrexcid93U9KOguteRX9uWt3HqQxL6QqUGmyXgix7KKiD
IE5dO6r9SyjxmSmi1M0z2cqsBQxQvnRDYZRs1HY3GnMmYMQneAovS49timqGCH6+XUhKxtmD5qd0
m3a779MvMyn+OpF/T6klUdvRcfBwPdCchGGL8jYrsuXSjyq8YcaBEl1dYzC7GjXfYzqkVax+Mz0U
X/TJz4H6ZUPmc0h7tpGhP/vEUFWSopAT6NIYocO2wEjaVJ39EaYgsVmsGlVIjjhN1SGBk11ILE31
fsKYa2xQf+Wje6rbQhYk+JAUFc5B3oesP6iD5n6SR2oQDVuecEh+yng2LyB5//Lg/xg23inFSq9b
zCGZaSYxKNBvXPW2IeYbumvC6qKMKeC6sYxklEDJjhT4txKXeqi875S/3qAtjM3ylaZkbvsgtLOR
/cgDjpbD40paY9/X7KsK1l0XjJmdUtSKIP9W3JD/xJlulFc2b6zAXADBjgrry2JVOVVV/SK0AceL
CJvafrCekPVdr12NW8ewjjBt3dI8kLS5+VEaH0XXT2WIb8vda4oiprM1DVPQADtQDFVwLl0WDrD4
bCRz4Elmy+yqskuWtj8YEBLRhJFKiPp++sIXR/qIuOOcjjKeO4Db27B/Drb0K19vvFajNbN6uSLZ
KGdDD4A+e1mxqaTTT2aE1300JxT+LNXE24aiVwcvslqbV3Cv0l/OUpTrHDjTEOgyRaLoklqaIjtD
OJYrPvLjxOYkYpUa/cqoeGRnR2p3JzOCLioSgifpfcJrV7rdPxVYwqBdVDf88e2vlk83jjZZnnwj
bhSfjhDl8nqVbNRiMP6qGQWdqjFp0pYGlwv/HLz47UhY/7yTIrXhp8z9BSIr7dZjJxRQIYV4tBPw
p+WIbagS3ddkBujIlkQbEM1z4lQDU+JCTd222gnG1MadeusH+I2SksoywrdTLTe4sfCq3WQO1Cum
9iVfyymdRllugZK2+VBbsSSS6j4KtnJ9xkZAKXJVhjC/Etdv446xIpb0sfL4Ci9y7zAA6GdVm1fU
9ni2XioQVaTsF4jvpTza1pUjvtVJerMVNHwc7u93j0Dk8RXD4YS5hG/+OV7Tgb0yf9WDnKVw5wu7
CDT8eWRmwTXX/BYH1nzAdsbHn+zCvJNwCKzWec4q4rnzRmeidDq0xu2xu3is0us1K4I5kTLv+Lfp
FcNLq5uKHr4WQ/XIK0GrYrS+I4OHwJFUMn3EMPhGyPKmRuxIpW7hSKdd0h4keQDQb6OTxbd5agBH
wiOc/wY7rPaAKiDU0/HyqnnChF0RYWMSGfz4mtPjPG+mqhscnCxZyqlIjiehnrO0nFQzX6UxR12D
OQv5owFKoi6UUDkGM9frwSK/oSCXVqCMyH0kioTUb+OURNIVWdvr000Svk4ciucUBSxlXd47WUXA
/EoikCpqY/Ni06miDbuhh3SQtVR85o2Msf+yxUbMZroRnU8Bxb6/8ZoexDDphlIAqWWp7gruGuGb
U58NAeY5g5v2ViiQTddBnNvnjCfkJg0+o8f3ZYzj/DGZIQ4pixZz/7TRWQ2ZgLhBIu4ndzGbQniz
MIQScEKXc5T5EdlqfPt5yVkS7uu4HPWrJIvhhLRjpr15YKAMznUtctEOL019CMWKAV/Ab18sY3hA
0aLH20wJDH/Sr9m+EFtuPW/sVHTqfyKPGX0dHMM9+CmYrT5GeeI6k9QlkWBpm5qyaXX2fbzEUiVy
eMFYNjz62yMZiZP9GgKZcedlFGfESHHjdqKMTghHP5RsuJOr9Z3kJhep1uD9fJdDAJ8X8ZXkx89E
UFFrSb63+dhvXjDmAh9Ab/KyJ9iqpCVPxPK2QiycExo89VYcRaLDe/MnOOyRNfd652wYH/yLjGCj
rbZWqz+6lgPI3mMeYSX74yxCnJ5WkrcIARgBly+LucFryhLjolc0AyWfvUv756cj3kNYlQyHcWiK
uLStega/+yQG1yVjuAQm+/Qk3KucW4RWUyey7dh988BHeIRU2eLLuIVpbxCu9zXJGpFOoC+3P0BB
T6Q1ZdY+ldcrFCd8847/GL7gUt9qOr3pqifIprilG+JnjCeRDuPwEMPBzHuyUmQlp9UcJw5ilyCP
jzB/THmMoYl5hp7jccgW6g2CQ//CcFXCrzqu/dx53VVF9/WmfsINyb8t0qLrZ2jgTnhJsFnv+ZoE
KmA5ILxEz/f/1fGKoOaAIVyooQSyzMXkoDt5096Cpb1VsRXWYX3hUwyyFBI/aZGy6sg+/VKtno0m
DFq4t4vPgxhZ7ZesceMKc2gpSd/mekJ+GuUVf3GG+x6LazslNnhoV+64KEXNn7Ythgg10Ezzp4Jy
D3HC4UIZEBDBfMFsIMNEHjos8nVBGUg6wWqfed6F7DC35P4uVeYNtz67GdT3INIzbwyES5o4WJYw
XwBLL2y2qqpxWFP+gjsp2DzVTVIdUJjPSoAAA+cVX2MQ0bc+uSqTNR1Ne4Zojv8n3r59wm8l9OzT
4/RP+fmejEgdoJ4LX/W955hXGtQeIn8N3DklR8o02FGiP13z+ymrhtBQSPPNA538p9B/Vvs1ihui
kfQOfx0x+WXq3Xa6u0wfZv2K2+vAg43UIAP61XWDb5UzW52D4ab535ZtYnEzXb08Rr2LtSQQfO1d
1CjuE6Nf5VEpZdozK7cY6oEq8H4Wb293emEXT56m+c6QMLXSsRmg22M9RbjRjfIFSFN9NGKK4Dnb
mTAMwth3jgYqhZGGaSPn0lr3Lo2G0rWXv3n7+EfCge++Lh3TmUT4SWk5oQ1O2fv6uXlQtWlTwJkQ
EKQxxLZhN2npb7XYgIfblRHKol5Y+rv+ZcgtlWNM8hxKQKdmr68yhRU4gySey4Q1nVmrreRzWUH5
yq4slFcjIgTTqvdzgSNq+229B0aHPSqw9CzwpAAwcehrWa1vrhcE3sDo1NyDE+C2imTlw4n2Kr/+
bPf/9sd1uXG0fRN7zpi/bl2m4d+9kn63DC42jAul3GK7WJw8yYWKy2veTZFY3J0K/OR54N2WOwLd
McD6cwTEbNaiqfRamd/gELHH6Bk89oEKL3mFp2dMnhhR5/WA/UFi8qA9KYVnEzZb0VIspaXEHphm
W3e/mTVaYoY0nmmGXudGuFqnzC7aEr3LZJstjCNu5EZNOglxKlrCliIiC55VKGzpVrmLM6q4KyYB
+dJ7NJClMoMfb+e3pnzc1Bje7AsYZYIWw/vLdt02BpGI67TYHrIUmfMYCDZpbKTJdWVtbDgTmYvP
JaehrNjU5Gbdd/i6TW5XLCIEtG+mkbZIHDI1gAGXsn6dLmY9ObMHm1NUZzCE0IPziXO1bDfivyH8
RxZOMc02ipsnr+6dTJRXKY7BgLPYRfyaPXaUTDt/CCzA3OdRbpgin1ts1Lna5UDmYgKkyu+9LK/o
aSqb4EyV4PqjHtWOYndvOErGlKraqKBv1dRSBZQNcglwKdHI8sMgRMkaOoZHfYtmv1YD38lWs1mx
rx2jb3jtEAWBd8jhPyr+pgcMq54zkefkRF3ZE6Sr3OhC97DpztBjeOpi3g8jN1mNa0qMNu0yLA2N
dm+X/rJPJ2uc7IGeKgMX0LGMLvhRXn7iEMcAabOX5kJRcUjX1XSOtuwwIjlRlr6gi3QhztbvRTOY
WFHjNeoE3lSiDz/6IsxA1XWx4qnj/12cu8EaQ0a7CJ0FOZPExRi0x3E1SAFChdWjTtIjANJwYTW5
R/LJreF3eT2jpNaYplbHSTKl2/tDDgEP4NPqS6mAR4qfwK51Iar2R/KbqjXIXuhVqoK+1KK5PnmE
5rAjYK8KAXcRC5tz0Xjui6MwOossSBGTLEnmi/zc4B/24f8bYRgiua+AIX3S2IDiYk8MdIkRaBKd
miSIQcWu4OurF09Xi4THGI711Z2UN72HlQoHAE2n6OnbWkc6cdbqW9GkJqzP3uJJwjPX10CynF9j
vsyIOPJu5KgDhArVn1YGNwNNu0KsAdvGZ8GoyP/LdjpPLIv6CUNeuSrwml5w1V+iefQ7Eww+8euo
lLfg6QRONynJl8u9Z360DRxy5duqu1WnEewuy9PgNu6qriAj6Nhsjaxqe7OzKpcGmnMgvDs6NooY
52dj/TCvwNatFMKeXW+zN9yEo5y+0obai7jOQmaVCthP0MItyJoR6ZHckLwsXHsxltEs8EQI7/Fj
EYoNrurcHBBUr5ftWgXDgfbKoj5r7MfA6wSXiucUHPd8S1F4qiPLi/V+IMhdFOnOCSjtfzNi196h
kLKzQPHLOC9454icfy3ofuXm28g9FFR9TjIamx30/ZjoPAhtc7aefMy/bMjtUZRBvtof2hhNB786
l1Sv6Yv6DRadRWtGXTH9YWFVWM+UfNXERSFvf0kq4ubUajc/4Liq8pjK4sxT04UvpGYFXg2s26Xc
SLRFNBLXxSsoKyOUmNBqCxv9w/riXu+nJ+Ij9ajMW8MOmVzclwvtzBu8jpdreIS8a9H9VKTnXhsb
lJ325wP1vRzScTaNc4qZFc9LhwQzxYVQ5rNmHyd35T8vlANJ+T9vIx2tHBTz1tC7ec50kvjzZSUv
VgK9S9n1D+rAyqgBiuzKgnTFg2OEKROrEE3dtyObkkgr7oFaNouqr7FEP5WyRbMs/3cJHB9FGSSQ
N6ToYQ2cLVMzSWrOZ3Uptik0lkf5qkChTzOcefCssorzWimaaPLvX9K6C1WXOE60gr23qObj3UYH
rLtLYxnlSVXIqQG3sCOsss6pjnmx9EVyd//Ve9BUSefHmuuqSv7v1n4a/K58oBcACpx0Wl4B4l3x
yfBlzRxmjMiNoDykHxDIi0mFXDnlPXDV1s4jhjzM1cdg+nFN+DCXWSyW71v+Icv6oAlyUBLw7a/c
7n1SfdRX9LJrE2JAa4rOmG8oSdNu3Wl22V2Fv1ie2LIq3Kxt2gyb9Qq8G8an9/uk4duERijEo2EZ
6stbWQROZVu72oyAiufopXja/4+85xDE0wPaavrMx3xdUc82Ixu7uz759r/LK9AuIbobbSr39raW
uLSYIFck/SaqictQ1RNgIWKUvo1GGn9S+eRUWk0jlLEeISxLkERzCtldQPMiGWmVzYeQeZdFHz9M
vjkXN6fReAmYTsvnIy2KS60p0d+FuO3oFn4JMLM+k6WUp2tfQB5jQc5p3mKmAy+A9DyWUhXO6d0Z
SYmbFoI3VUMLNqL5XpuLLi4T5DOCiYs2/gDKDvMPm4kWDIWybXqitLnMDNLakwuvJshBoiiM9mgN
7Z+eNuBzQx0hfL3nQ/NZ42eZecJAlB8dsGLA4xhM1Y8RtLM2LeMWbeSBAczSaycbkwd2W/ie8LUi
WROZlhyewqYmomrzQiHsoNFx5DWUoe6JSu3uHx0u3vknSKWnKQPILnlkDb97Er2AF5H0dihwsps5
2Smk17wgpo61s1NqGvt7v8qtQfdf2tSoesp4l0lPV3SvZ2jyS7uh5OGrJWTwJX46qcl63ZM05Xc3
jgXCEin8GWYHq2KvJF4riADIi8RWdhhDq1gTSWPsQlOlmbxLHER+diuGN6Uk2Z6fD38vZrUmB860
qjC//k9SfWMGbXmOLwH37dRHZhiMSqeR9jb6Ae3L8SG2cfjGdbQ52XgN3CJXT+4vqG6nlwnNrPU2
zYfaOVDk16A9fZcrEFgA6Pc2stBqjdsU/JUQ7vQ2ZHTvGfE+7UIJdRT81pctaxzSsNT0pKx+6gJz
y0ekJJbXqwALeHxNO4L2QXbfAao9VsXXc1BYQ0ifZCqkvSGDpHeAzZwXiKUwPY+cGV+GO1YWzb5q
SgsGplee4pXlLRotJBwfDtz+geRf/ozZJq4YXDOibLitXkWzEGiIYPGGn84c8nxheC95zzUduYgC
A5/pZFlH2exjgXQN0q81Dj1fndxeb8QBpHC/Ranme4/Akai3h0afpeoCOBl45TpiYkHcHLVHQe9p
aCEfeaqhokkbM+Xuz/l0CbZxQNcq2A6h1jFmXioKcVQUZ+8YxA/nU0MalcG82/CV+6+ZJ9ojprRt
cv1rANEOn+9vJmvffIVeQhiHsfBc0N8XqdVGkUJK5pKYWHz6NG0bgY6vCs0ydrhE2qFya+Xt7BE2
FSpSOFWqkl4cpVfBX8HRxu0+fgkgZk3NhBLS5M77CJ5sttEvkfqBgMCKTHAYk335AgV3VDj8RVD9
XKcA8GhVUSjr5RxHHWwH3JBRDt69KG44uyr0QbqEVAZU9hybm4/vv0CjWBxfALHx8ILC8Xv2l3IP
bElsWHdZKSZhSrGdfEIyt5QFtErP0B5BP+8YSfrqlGittDdzyEdO5A6DwaWnOyv24OI0QY7mP5Ya
8ljbu+XlpNDF0Mh42ekxvFdMW2cn40jq5e/TsDSdFlDfkT0Qi8BDwENOmgJTYQlYRDpz5CU9ClW0
gI/bK+1pJXo7qCq5/kMKYnyUSZ3K6kIcCfokScj8m6zKcOde2eo2hn3a0t8jvnQe6QkHgMRDGMlT
kvIC8CYL5zsBeiXzEOsiiUmtGVqFeLuOpZMPgVohvDjAJJxgbFD6TAglGSbmipizwOonpEMwxebC
nBC7MBzWGoLPjetSWYqBgMZB/48t9sFJBhWP5DB+lz4uV5LPlBOYTGBCgaS631fu8ceTzIgvfDQH
bw7wCIOKI6th0yiULy3Fr4KkkNl8E2oat4aR6NDzU5O83wwZV5YuRx6Bgj/KjdQzOUzDBWc2yp03
/YDgTBlGVDQP9kgPu1s0YwORqm56/AP6XZWJeJANWPuJjBDTj1gGPReQNgpYlej/rxtYcyWY2+sw
SG0P1fi2eD7ceweWtLiL1DDOrNF9x4bry8g6+jxu5pnLWS76FDlaC6mvje/O5QbXjqzo6xK2xsLl
Ch6sggfL7ldQXbqh5vLLJ6T+Ll7QqvlbW0+a994soq+bdTyHMircQF8+RHQgWJKar2yBODG7VAz/
9XfE2mUfxHu97PtmsSEflBSn7eAJIurtsk4+TybX8YWw6vcLW0TONQZ0YtAfyuiFgOKBcp88/Mbi
ECtIiyjxI0eh44e0mletKyUHEGPbyofgeJUAmZYVx6DgO8IVIWCBw1IHWX5s/oIb+48gMsViwjKn
PAkre4EjX3ViRj/TKe9MXx6ml1KVniTUJ4hIGVAs+l0uqZ0G9RUxP8G51KgkyEruzoNjyzh5OCBb
CQCv3tnkCW5lNNZVO9Tjh6d7xAYp8URrwoBH89tcO2RF7VinysHS3s1zj+MnkQd+n2s/quKdHyG7
H63dYjnQJ7bsi1ONmgeMq6w6CrjoTcC6vYUFuCgDnbY04bB06cH1opd6Y/Xd5XfyXP3n4UOyDj/I
NQcj0DhdCgLac6PP03demGYGD0OBSvarBqtT4AidZGhkHfQhYx6NHWJd9usWx5VZG9GC/6Y0Gax8
xcGGAahGKBcrdsnx4pqHfUp711BE7C2UMeZm5wZaEp6k7LZzlgY2jfmrW5r2RdFHRmxcNWmJfyXJ
z6d2iAdXedsp1lSL8vD2dsawrec/6705LgvIZ5J9TIhfFo/kSPAar0s4uOh7X7xd3ytJmIQSucKj
mwUbuZtpoUciavtfS8nOFaM7V1rcMyQ06os4rgLXi6INlJuRNTMpJ1pCInCoAEAV3/ObMLw1RTUC
OqetD4T4O5HEwR6vs6yKBJaKDHGkUeGkJcIpiSKzZyFGZlAxU6t7zH4GkSlGeq6q32nyC26wnBc/
1NW5yvq/mT1E7AO5RPYSgQ3pX7ir391O4NIAWSLRTkZDqCkS1QupBCuqi9yR4UctZfDQeFoZAp8j
AT5jODfanAL7eDezpxOZHYo4MKolxlah+EuztBugzT2tOWPODcWqY7vlPbO7/OG9oAiO3Gb8ryc/
wNneBj414W3cHV++rQa8CWjGOfUrkSgUkMY8Z5bC5oG0sBubBhe6SytObzqhTuS6TiqiM3Lc91py
G4hqa8MrRncFR6xQyeTg94Xy+nhlHUeZTtumTadufe1WVlaxAeZGUazdQdSfDbKipq0EySew8tlW
R79Qtdvg2zBJRToSD7wYOJkV547QS6oYkfRoWaKN1pBiNAMxnLDHB8FPS2QHjji1xGXeIjmCNRNV
FpIP7NWK9lELe7i3JTQ1SIkl3ZNdglpATKc6OmSx8tgWnJfPOgGbQ78aarWV7NO0HLBhCToYdO1X
rhY9VFuE3AZQr0ZJg1rY191o8YvPa2yQY4hC7pingHwmeXd+0N96sKxTEF7/Fca6yjWcBoWtnheN
ONkwyOxq650S+NxIkvY/E3hAv7gZq9KEq0BELtr1+AIhEMrskG7TWHB7izpY3FgdVBNvNuIWJ8p/
uzTIPTRdidH8OQkoXZ5yT/nPbyHJlLwJ8j4hlNmF5mg3AKZGQoz+s6wXQCigvh9enS9+PpIfPw6B
KrcgPQ9uTNXb/vgCE8zDCsrcpnK3H3MghDPbcfP7T1KeFfJlwGU/GEaIUur+3Wy34Ys278E6I4un
RIRUIUW5x3DXWV9GKD6LstUPi8PUYZ08ylvr2tJ7FM1YivnD5jYULzfcxYG5pEKynmiJoJv0knDw
twgkJU3R/XjisrT/irNmem2o2XjsDGrOyYfZhyCl9HmfgtDiyDE3rbHtDmy3UhyG+jDuo4h5krhA
e1Of+jNs0J6y+B+fNle+/KeozrUGz2ak2nv19wlHu56iiZZCggFsHL4GBgBd3cJVh4lDsqQt6j59
sI1fpdZcZvz4C3rLhNoIMXxywNz9BjZ9stXu4uOXj1VmQ3/+ILI8t/6q1tmgN9+qupcEWbTYp1e9
xczlzsynfBjEG+D6F3b6Lol1yaL4lZ88h9Jz5VnglrQSPyKFJo7Q36s9/Ice+BmktukiG6WxtrPi
vYbGe3Tf53m5x6IXIjt3rketHi1/1oChPQweLN47kU1kHOoUFYKTAOZeeh/WKRIyGXbjhiyHIUJ1
2luramLYEfkrCvxHUzH2tuoy0tAl+2NipXJbJA08DFTgxvh2rDOY64XvzQfWh1/EoKbIkwhQNILw
lIT2clOEFsCNMyPFEelyoMSbu7amnPdCj/9PNPKZuIAQ6iDiP4kYdEhoQ4nSVketmA97OhzvM11q
9NBgaNGBUdd8OiQdLZ2ORfLx3ZOidRBdk1FeoHMtDt5hWn82ACgcxHJ3Ovpyl5PM3jz0/wH/wTDx
pW7TNdYybmE1cNT/AJ7tvRHac4PkT8pW4kUkJjxlH75hxuoqVxmWNFjZeaWZKusDaG2oyzHlVT8U
1OEmZSDGn1tPIMKwLwhPgMSbGE69HfOWsNj2Tf/TDk4d/cG3vL8ZJTnUwsI/gVNIIRgTo3TL4oWY
ifMBjJ07KwhwrQEw1YbhERGiRT9o7Daux4Ih31pwi2w4UVwOvMPRuFDBNwGEkHWuoipF55vE0va5
+GKntwf0zvrnV0+kHl0yyXXUpu9u4u0Ew8Y+HhTO3sf9zIIQJHxEEeLMen8ePHgPg7cfTqV/PAxq
sViqGRJlygDZTGOZbDcb7aoQ3k0+6FNCzHtHbBZ9WFORk+h6BhVsT2yOn6uYBllyePIhlJT6XfiG
putKEnRNVinzgQ+F+4352D4q/VEioWZqJQO1qcr2hfq0LxVKAaLIW9xzj6ImyU3yWJEAtyxCWdQn
EEAVCy3W1fAR4yBHVBjDo5NdEaNatJcDC9ZNryEfitQw12PPq7iktcyWXTttMGZ22/2V8BODxhKo
8c94joJTg7JpCRQMGAGCalqKbn0+HkK1BSq4rNLD+1Bn6MVGkvhxuol0pXkq0cUAxtxOpOWb0ZUV
NQ3LE5jltFAuqacJsr8kuKCSgdZtDIvxgdDm68BoE0pj/EL/Xd3iyeRSN1pq51EvEwWclAy8iKww
hsdOSCzduR3sVfMqK6mE1oz3ZpkxKm+qJKKVZYSyKdXMZ9NGvPWvwf0mjSpoGBTtO/1w3HU6q0ev
UYYkGkdRD72cQnBth26mGYff3SMTsNd/1eDZA+M9C5j8Ehuy2/iM97rDOfHb2ENH+IZ3cEL5QyRX
m5fU6xpY2TET7Cs/XjWtVJsTEVo8zavVBlp8vp7AWju6Z/Are+teoPbRbJ/aJab4DV3wItjPD/eN
lLF2UwjrM0nLp/p73dPvV/Q/C3TYsNonAbrIikAkgg8190pc/3waIwvuqHotZszlbE+gBjPofsZu
oV0ABNscwkMDi0LzSzlegdjs7BpEcyyQAYJQPzF3/YZu92XclE2y/k2ekSYPxwoJ/PSY3BEYhLyy
ezb7c4A8abGASt5Wf5V1hF/QRTg7+lgQcV53whfKb1vmzkyy+Xjn8AB74Xvvz+69vEfrRnLr3kb2
MkK656TbPi6ntrZTLqQaUF4RvknoA9yGoMqk+pVRf4rmejjZ9P5A7Dm4u1+zJPE13m3OvXJBdqix
kX/oYl6hDHlmFsLJAKFFg1JOo4qTKmeqv1iUr7M5lSPD0RSGE7hAgTRpxOvmqrdNhBhv+SHAPGxW
45BLJL8H/YNiqG8ZpuZDFmV8EqN96ZmQHnCrRX+TIveDwPHCoPbwQQ8FdNjlzEbyrkj2KWTuQoZp
peeDJcEyjYxXI3GQixQuaxRqavNfxdfh3YFwuJs1exWOyvYqJVzL9Fsw2t9wgvdhnOsPHhR7AUeQ
fLWRJy0S5cbuef45DOwTvvv+L2bHrzX2mAY5Hi8dLlr6vlIxaAHsW8KWHyFV5KrXNUyeqeznYELp
pGJvNCpMM/kbHMVCKdmb7sSeOVBQtJf1oxTr87fz6auoCTTi5u9o51k8fcwzAqnMw4lVsCvIiOdM
XGv1K9Yj9+zfwSHK0BhXotvZpTgrJUwh0JRvZs5pBU49IplK8a3pzbjtYwL2Sx5g3whraNZi96wW
6Oii1CPH4IAUPB5SLqXn/ftE3c36pJD558JgwOQIvSa3PAF4L5cAyH1aA9gY3YxX7sBYJFLuZeU+
IWD7sxZh23iubHuMjtfYO9y2CTaC2x3wfYJf7PZG9yUmhT2J0lXsFPSBnUGypFEbwfBP0BAKMk54
C+EGWxPBulo1pGRG9/FHjeqydCGwTCmehSBN7e0kZGbKae+2PkJBPa5BAkvW8Y4A+O2rgsBlnuq3
HoXt0CwZFKNVvUofWmcli5dCrj6V73Q/LKMd72lV4ADuba47Fneey9EyDG+GvRdQPTP4+QMXbdS8
GbMbYEpIXbS+JzYRgtrNWN38u+eGKPH2meYJUEsN+whvJ0B6eM73HPobfPc3ClTJLvPWNU0NOVae
hqNfmywuzcyfLJsHbLgpmDflQY4k/9NSAwlmUINOoa5baaCcv7QKvroHHb4kU3jFse8duIAJtWeo
O9orCjl+EkAnw6cc7aBUjnmBVlZPrTOIY4KyfvFjK902l0hJb8UgWALrN9kxL1JPpAazUD7jWfOY
MTlRSlS33Sm4kkG1Qof2xpR7BI0aH/TBO562F2+badrMp3CvbYzDQv4UAtEX5+o7+/7ppLRmsF1w
Vk7eIjT00HM2BxF/A0qNG9tGCaa14YDyZsGUCe3oAwANShB5+T50lDK8/VaYAANC8dlMl6T5ddHN
XbzFdWEnNgmpshnpHU3ZeW25UytVoDNmh3PqAQPCgMEW9p+QkZ1j/raK8YmdrIJJgIo3ScjMWSw1
9MI+sZl28Wsh0tpI8RGDPyhWZm2NmmknqANhsSQ+if5Qn+BPFR+djeWpObFzQ7lbJpncCEm+giKr
5qcmBCFu7Vy30MgY0iZA+EwAZRt7t/1Oqi/adE3YabLsoQX9HpBuXbXubQM/04QKo21MsUdn7C8/
urR86M3LiAuj0VNHMxQ6XT7pctw9L6ekSDasFAVMvMxZqE6QknuPsDc+f/evsQGaCgUmePQZStBk
xacWeOhKdXGB96lPnAAbKUXt8x4HVmRT006fdROU6vvFUyt+hTH4iEUDojXtUE9Azw028umiYcAv
CwA0XngJoDqOd0baRwotxGPxMNpsG/SJvl1ULg/kgCYihC64NjWKctvz7vAj6QnKCLgR59auUAuR
rdBnFRbL+f6z7jBtw7g3xdT7vgkiz//BoHjnf7J+sC5AeREYOgH4dNhFzoWHlMTrrdkjRwvR9yrg
BB1Jy/HVVRQlXN7YEisb9a+GaVs4SjeWfUBuWpfg4eZyVcGfDlgk+bqNqu45IgnrP2Nj7dHHNL08
AMh5a1hjDSY84hcsH3I1FiudfKEt/K+j1S/Ja7Koe7QejzmBT6NCrmqaSZDDyO/7QbwCgdFqQ2an
SqyrdXVfuYu+kuLBPCNXiRWZgJmSZral+4moOlt5fM5XiUr5aKN/NhKnFdtdD/CyRJALtVIcH1O/
ezwej7zUcSrynzKD0aQDJ0xOADeX47IJfH9L7IuV/xeT2PiejpH7uuIm7YOHoEOl1vHUSSw+XVD7
0mRs1eleqtRvG7+w2I1SJgWA2gPv6s9r8sX5dEg7r2KlgmVB7dMhde1zopLxeR6zuBMV59SUyMb0
9rb44l9kT/pEDb2Evv0GusimHPQakCY41yAu92xth9SPRumOqqqnsOE8pKk8sHg5JcEOq9JLH0wv
XbAT6WURHaqx9OfOEuFCalE2zNxfbnnyPGKsK9K6dvZ56q+OIXWfkfpZSgmDEorRuf8Zk/53AlnV
BhlEVn0iHSGOHXifGKX43UaHGR9SlqtZyDFII+MbMfP0TiQlU1M6ZI3XxnoSreXqRh7LNeLQDgFW
4Lm1RhnK4JrjevjiwgFcJkW5lfCZmdsFZ41nGRjivb0RpCqYyVbIz3FynF/4zxNKjL5XffU3QgpD
uN6BrKMdsgvSbdKjMJkXTV/AJT+nOnDrgKS4bmI9u9FxQdtIilwoC716hZHUDzm2Fnkhf52MsYRJ
jD82lnC0q0Ufbe4urL/pkGqn4GxsyjtZ8TSph7mt5YksjlFZ2/yJJ9C+QrhK9Q77+VprU6udrTM4
FGSnulCh73rDiQcsLhULx+HD+ZMh2icA7w6Kgf9neMWFNXneOrjeCea5LjnPrVfh1TV9DLv9OzzI
fI0cmO081/YyOuArUEHz4MGag8U7GqsM6OVVdTZOMmY8OWwShPdobD2cKig1XLVhXA9EQf/ncK/c
Y/nqHlcWnvJuD2amLGsdphwUyEXNcBrzdARmSiWwnGf+OVwCBNyLmGXCkN9OtQ8iZYRn2JWYRhdc
tQjns27TxiVeTTEkDld9rbS8dfHLGsONLrgjsm0cFT2aTd3kxqqwBhQiIoL7m+oLph6iEkCm3q3a
OM7cmbMyHo9Bnj9WuGP0ye1O0QRQQ1hqXyd6vHv1DfdiBxcloOrx+lv6ikhnd0TI4IpJ9fb7/AQH
nOeM/ZQcp5zVBZg/CjbjzHHzzCxvRwgH38GJdbGks4o0Q+7+uqniktC/O84PNJqhRWW3TOp8c+vb
fDlZ840JOIUmROeYAYiqH4RsKZLgwGCMMRxIFn8apu3Fx0i8cXq6ffrh7z5XnJl7KxAI/IrLfqb9
bLHPj08T9CfvEx6f1oTAxOfb6Or8670dtT0Bz+tc5N3xW/fAmpqyR6+U0dPVa3scuA7cOfzDWJzj
4U0vg/+4rqtZDxB1TKj400QhosfJPplrKphvYYzCyTO6IFs+lCXvPni8Pnrdq+SKe9uEI5voYuOK
Kh0fwBez2jt2p60Xdcm+ahbZJ0mcUoS62tyg4tKTpwhWTiALs8ZxbGPdJ/m5qy8hvyFDiVfestbd
4W2Sp1jCgBVTvqq+/IKzf2ExPN9z0RpKbcCwc3/cIR17tC30sVBfIRSGNs2qJ2mXOPlnpnmilrZ4
G/2KNKf22U49FgZvUh7HwEGCZnIT+uUoVpz+cGr8oN1lJ00G88Mz0UrcNO5EZ7/FXrNlMD/lHPbC
fE2q1a4oyMJo8grK0V0hY/hK6Z5vNN13RhzAtFut/aO5Yq4Tltu5bj06guhpK50OtAj/pjHEgDgW
SYHFqTm9ZHMb4bHawsks2ckOaEpmIlIf40eHdz0OOxt/EnqKV5YOCf3E+V8uqWopDayfSyT7xlKa
ulJuNRL/HZ8XHl/Q5XS4NjB4cvIp7cuaXccr0vr1+lV4MB6Gw96YmZpthq/F0XgvMwD3wu6NBggn
P3ZqNS3L3ZS9AgW7+dUFGpUd/1sWpdW6mjDIBOsLYkvwLzWa1l+l//oAG/vbhKoCbgUU5szONgl1
SuR16KaAgWJMs8E8gXoOq23iXY4dxaizRk76+ovMrFlkgADnQnaiY65S9nXehqcyLXpW6kYDA4HN
xwVKM6XzjREaaD1Xf/xMZnbfHH8I/EHBCvqwQX5h6xJMgjrJpbamrA+QFQuFE+BW+fugaop+EDbo
mLUfqUfbA2e9ry43218FMy7phtKK/mCvlhFBuA0rJm2CIbJwu3GvcXYoAS7egcvg/flYS3GmKBXi
wkV98uEDJDOOwjoqJXEYE2uiH6FbVaEzDKdnpdEAf6JVbwAOR5Z6RdOzhoZ7rFs8Iub4Lmc6Lgkk
ISz/2Giynd+cQKiC/2zUdKYc/thCdM52qs9X4EcCbv6ak0uTac6UKDJobj1VGyX3QJDNjkCc8Ild
lKIKppAwTAFn5hVpk3zpvKlgau+AVMT2ssfhjb7n8c9D0m2/Tra0b8ugbmrBtofyLy4qG4EkqyDB
t2/n57CXIfAZeo0k5z06q57+CJUmGrIs7rKcbM3zBY8coLesSlim7Wyu5+4eKUTa2qk5CtqDDZSF
jqqRR5xG+xao8f53FmGVnjk3R6uOrik1vYRVI8Fg65Gy8QhTZl3y4fJV6qHWTo5aZZNR6zsMLweY
3SwZUND++JEijwA5441OzoRHYsJjvNQ3zg6TnYvR3ZK17cdUFp3LakACE/5ExwJghxUuLNXwXpRe
u1FdVpxx9PZPePtvfao+Au2jA3X6/pP2nsnFKdQzYK8jZqmfTDM10VjHCbqEavNSHSmm7Pr2R9Ay
EqnF/YKEnbaKRi3V2YGkelgy58EBjWo0+WTyaSqljbk+6JBlc6Gm5JlWjcRBqUGr0q54239vbny5
Q8HepPqlRTla+m465DWEw4we7S0G4Kqv3NiMJQuOySpH30UzPxoRISe8F/UGia8KsGo3P3HRXc5O
KrtJda8z90StyZDeWLUyCdvzO1f3DSAbrunWOIxnqL776CIDgr79w3O+4Az++YmC8w0kDpgGKMnU
dAr1NqJHSqMRbcAHK3fcj4jKnujC6L3x5HSmchGSzZW87SuFMXh0nuu5RllGBnPReMZMAUUnq9cn
5UEEpQihwsxYmnzmNLoD2CAidLt75VnOeA3rUHTTzgw8EuLLiAn7DpdAthNLhWyO75/oNN/ptKCA
E8rEoq0LDDWlqycDqKIDcWkSv5T1EOtHqo4OrrMmPWJZLEz2xGyDsWAjLFobhU8Wo9FVTVts/Wi3
gZW+TLxN4b6JxRQRm1nhWBIekB+a7Zrm5bLVuYqWved4fN4qsvH/0SVKHf8Q4vTkAY66rAC/ECfw
i4R4lzDnGvnAFvlf49BH5YgZH+ymzwz5pg4h6AFNw2/a885Tl6sNEFhd2PXrMhbUF/wMRT1ik383
wZDX+MbEw7W0cIasyZduvcdrIPNneTK2/oC2dZJXLSW8+MQ5G2ok4p4IvK5DMg0qxkENUazEtR6/
/1ebzsZPkAjP8IX+tfun8TztRUvEmmYDMG4rFPiO1iyyW5cUoTlwI+jvfTHbdwTtFfY3MSSHt3OM
+hqmvywBVNbYyu3WCtgTLu4ONuHNBFdrPKeS2wd0/WCW5bYxf9xi/kUO5ECJYcG4e7T5Z6xwF0+1
6wiRqfNl6WDUQYZr9aNJ6CLIkzS5Sdzy6Rt6nKlquvP5nRoEON9PETfXfwIerQX6JNEHb01fAwku
tHpQbZHBFHNcp1bEOhOT3Cq9ilQBM+8/+goBg6riHnhPqWX2WtD8d6cIPxc7ZUMiWPW8exSSw1An
zm4gddI1L5ZQVo39Ls+tdDNQKiMBoUgaynOcudNQuHMbTsuJ2bVMHkK5V+d//e+1SqKOoK1Cajr0
lK5cAstKble4Z+apq8yy++XbL1TNFwhzULquQ1xAkN8+l00XqgF1TTo7bZd5XW8cGSrCUbSZ69op
EelfrO2ZXm/bz64gEnQi+Ph4iY4hsp/3mn7tC82EWlrg8grz0a89iPqa53bno8Wgh9kQ0UEN5S7L
JhOx1K2/wsooe1sr3T3xgCTW0kd6OjPlj8FO4PrDgTU7Q1qK2IlT4jZW2nNTUfDwhor0ZvK3Oq5T
nYeo6mmURoqI7jhY2tLJIqXU+3rCkbRQMg+oYPSZ8bByxfxUyYfO5pI7y4G9teAIsWnxyjGxAJvV
/T5KrnZRwsTMK+Ac506TgzmVF/aavmOyjqYngmZbM1BRKs18CiZwXiEM8NntymR+ZdeBxjInaB/c
ormHoGd4W9j2tHTgQexDJhmItU9pQxmy7qM7goDZbW1c1j3lVdvma40rqB2DptYN6lafoNEcyZoL
EFjea16wp/dUHf12UPEFFBAdhCy8YJpqjGbSva07gsWomF+lrGB9x4hU/448P/aEKtCANlyy+HwY
+xlfqoMoOrtgdY6wPoU0KBxmEZEwA3wZ/4F6ELf02SpVmuXzh20gqhY02qUbjTtnOLBZln8yxSCj
r9cScMO+YD8dcLvCPO5hemDY+NovIJWKxwlSMGZVJqoSgLXm2dfctVDdQjlGxY/z8Dtick0EMemD
STzp+9V1fRBddKJPwku9VGiM862TnYCbjm6YYV0Z9HEmNTGI+rogZrWbTk3bXDh9OFLZ+jYgo6Hp
TKidomD7AOFPxcUDs4EarPNjMPhInpQtgI8W+CvIKpL19UfpXABsN5xvnQ3AVnx1IGgMnXxYELh4
oFyHPk+8Qa7AqQjIPh6STPAMyM87Kr1lWrBtESHGdxCxcjvfknkWSu0LED0SN3BllTyAHg8RkzGI
oYzFguqrCdmwdPWW60TPkIQb4ukOoodDRHd6RHQmghYamo3ARj8aLb7iFXTI+MzJ26hdcTR1xd5B
G1wjvjXR3pNkNU65YY24D8Cx4eiSHi8hdV6cxixEGTKtXSXJeylIPXqZpuKlpZQdXUKANCkI2frU
NuYaqHxsiu/bhR7jzRSUL3jjTs44CQxScQBD66rnOqXc9dC6PKzcU9kEdroJPjKMKjsasU593p9Y
oDGBzOkjL0hHRNbbVQq48jvDkMbr/XbMjpnmJ7a1+Y7+NnVWRlFs2dgj3jGw0zHW1GG1KKoYsQDT
VIpCOoEbk6YgQOzzPv0LUaZHsX54ljvQBNLFsYcCoUfGOgG993oDPA8wlDNzZYLZEDvMmQvEsOCl
yb6Gl2urSUBoMMEbxAPTargoW0+VLDVkoPZksf3GSlgiFquBBib8+Qv7U5IXKaDtCxz6GIaed5OQ
zAQW2WHyWIQYBz9e1BgQH9Gw7NKYhFKicUwzVWl+/x004YE5rPlrHF+Y1wCnW1SFnA9d8s9keGvK
U+X0dg7DhZYlLQbWaP6EzwLustY2U3MdsEeGG7Vrxx//UEqtL1WaTR0eLgZye6bFycWr7olXRaRa
CG/mDv1/pjouwEB91KvGMuaS5bcvv/Ywz6Xpvkn2UVwFLjGXOZEsFvW+tpfbvccyUnc0gemliXSR
8kUThXTvAid23v2/TuEE2MN+ACTvcRsLOkufxHrKaXkrWBOrjo9InWLPxweqf3T6Hkp9OIz9jDYy
WSC3KWkwVrvjRX1UN/ogYf4EsrVpA/BC8zXgjcIpuL2WbLaVCvA0jlWaR7z2eehYmUXlQWEK04CX
fqbOkSw62hNYOx3HCCRhBSJ4irXMOktE7Aj3uUeNftupZjLiNf7HzEodI72dCvyfQACG5iSs2Ulk
etVD1CouUk/pTCXrejeYRLndySezSSBzUKlGkaNSXp76h/nv/DgD68P74xLjY+A5ftfWChKumj5J
OJAuGIkXhwV1TuH2L0qjE4f4rWUgG2Jp4zAYwXKIshmjEF5NFBwmaEfVPh9EhHle2UYmhzfMczUa
fQEF/vdx2Zl8J3fFt9ej/p3luGIZgBYhEYSwVIzgnlk7uIKYHkhwT9sjhiI+xFFgA/+i2xn2PmBK
KaEcEpczg/hSMkU1WEeiNOrhkWE0DR3+8YwZd4r5zO6l5Bhople67wzB6+YK8CpmQJMBJ1Bt83oo
YcF24ofrKjfy1VhYrzfWSIYzSf0814VgD77DODJPQLG4Cz3VqS3aTJWZy1rN/HfzSs1dq0XsLoxj
QbtlLEx1MkuBwNV90QRLt3wU3amrW2xe+4q2xQtJtgmFnGk2pqDE/n29nzxYph3qAlufmsCP9Hvs
sRR9m67QhgO/DAH9RQ6C6UQWTG4FGAwznYt4udb9WAZ9uIKyZ5Wzu0xCl9f6o/ifkpXoBMCkoBIY
gBk16kKlXF8fZyQ20k5Ae954eBngrjiSsPcnyyJgSU0rYEnjlTyKrXnlH9tIe/1XReQqA4/Z7FOp
rYbGxeolh2eFsbcV0UVbfdn59TI9U0WtyvOEAyQoaQdLxrlAb8B1BadNrm0Khf/MYNc3eodhiq5s
ewGsh18SETQwonpgGdVOYKZElg1OYKGz2WiFUoDnikbluWHeGsbnIWaqr+tZg6JJ4Bw3EZMie+OL
2M/eGsUTD0jTMAbLk2FFU/ihUokerPkGrU0AztmVb0Bs+B5JTcOqQZ74HvotGQqOAQNMSz6yPKEL
N96h80vjDyipPlAq3dT4Z298aYeLYsnXC2nhKPp6PCLPzf9YG5OfJTB+0kRwmqQNk/DZBTE+3FRS
3cYP3gx4EKYMuG/U4bVmbJCA+JT/xsG2Gnk26ebJO/OxqBAgFpMjgY6AOaGciMu1pGUr0A4zJMuj
WBrY4hXeyaOYEXTe2nKRMta2ErdrX7y9bLY2KG1Y8gyoCRnRxFGujwkvYjvTVJEhnEJ7xQgndZ0x
pxzxQHThjAtvIiEAwCTFOYBmD59GOZNPfpIy9jLrWsCjBc5vjCniuojGNmS+RlLJUdVa1KQ4zuG8
U8ir+L7OoEVLkZkqrkFI52N+qvW7W0J8VvLA2BKJWaUxTRxXvcLfwH687Qn51xvCbhGCoddXCKJp
W/Bs2crx4zYaV8hitVTFkiVTo/jeZWYm/LRoiYLrBIRp94LgvZ2knccuThXpX+wPGku/EYGlCB1w
2+OdrZDi2bGrz7rvLHTEEP2MndqiUnGpXZo9jEgkJlTDz4VUNP6lndxxWO2ueztHCO84EG0NLCBD
e9z7d7HEhDMpMGMPx/8wboFMlQ74iBlhHGOVzs1FicTNLiZQe0DjnbjUvoZWFDf2F+oOMA9WIuZp
aLEoVUYsHaOJWnA6bWZf+r8w2biT94qkMUG1YRsq6za+cFXuBpKgp+UX7rNXw6TgmS7lNyQerAau
XC6X9I0iL4x5l348bGTv+olXm9mfh7CcM4U4MnWLu8pwN+KHmD/cUXT6ZCIZ6oxXbmPSK71XTHlG
A3PFzT/4VkhBvwTk3MLLviHGI7gASVl+IqFdGnvoPhj19R2qrX8aTs/mvWiHzPQlaUcwJNALtJfJ
dBeY67IziA2flDaUvjghfJCzyj6iXsAz6e58hc4bW8CUTxXS0eUOmVOy1NwiHpLsSsIIiODnRnO2
4wIc+RcRx2CI1klnvjY8oTgoXIZ3VcALMUk+EiamAgyG0Wp34E2So0qhQ7bea31JyKCi+mCUstk2
gfU05vxIUWhX+I6CoddXzpGLpRV0mI3oVWHfbdxjHdow90zvkK07m8ZIzp1rRJNVY5GB+cvR18sZ
MHA6wmdpNfqIQMaKGELGM7mVy0fNgKRb6Xqx1XG0NK/Wme29RpP1RBRXI24oZ6K5y8rYtFwgX4UV
GeWjeFTOlnJYhMcjSmnKy0qOeYliQsbuI8CnaXKj/n70DsMwhFXrydj9NuTyusx+rgzbiZy+IgqY
+OiLVpHhy6EJHEhIgNEfl2s9itBFKkjT2t339FfUELkvN+EkVLLYwjhwDe7sQZileEfMX2NcbX2B
9fKPTS+8XsYbkNiXfaDqZopQZtysZ8abocruDZsU0qC8slHYJgwlEKshauIoc/6NUcHlxSalGYya
dAntVEbp8dTo2jKkmo3MEHCJ1bp5nSZp3lbU8MKTxgyKg1T7bw13ewrZDnBLkstYw7O5Th1mJZEt
BUZocJTHRc3zhbDDUmu9xwiC+2IHam11+spbgRfnsYbezHw3B1GbCkGr0jmq6vZ/RE4bBbOJHbv1
E6NPwRKLvzpb9EFMWfIXU667L2XN/LpQ+kXIoWvc2ZSbEUPEZK0tOoLf3sOclv5Wbo7JyV8HHSwk
NLpv5DjGnE2q+dEwBdBkfxCpOTc8xunQyfEhNI17swxRQirsITQL7sSua8Gkr7oz7fMmjakXHHDP
SUO+l/DLWdsnHc9kJSwjL5rowYnVDl1GxpBx8gdH1LU0o9ZWYCkl7NdROx8r52FAisDNLHuB8cyM
SRoBm+T41OMUSLZs5ar8kc+31L7LdUylpjj1gpV6JO5Zu2gL1bHoVdokip6xcSfxeuvl+bHdXdoo
ullGV6jdOS2Piogh1awsRdo02pcxeAS+muHApcl57WtjTNvZvPsqYdtfqQqrI07CC9e2jujGLL1R
o1rWvvY9BlVpQKDFN8H94HWZCmqkpu8uj2AJtPaSQ9DIj3gRYpxlAH/f8YbkT/RnS/a+0ps+/dHf
leieps4K/Xtfj6jquv09/wFhm7rbDYvY5c0M1ttZg1/jGVz5bcASM62a636HVeY9mqvczj7G0kQn
cYvT0Kqe33BGWpSnngTH7Rph0nb/Ei+c9R+7ICu1m8brbB4a2BUx7LD808EA3+Dd0doufkO/CPMN
MIj2cHGBc2+EEVYr74KUwDjVVZRQ5PLXH04iEOKMXYQKmiabDIUk5xx1ya2VmB07LNh9goq797Co
1YnM23ZvDx6LtD+/ZyQPw3pqFh9fS6/KdqZK7cAWD9siwCPbNxPfGYEVPgjOBc6CEgz38TBqGXx8
M54bRpjCE8nm8AimwPPHUaTNFkrwFrKsJgJOi2Zy9VfaCkD+GSfzGCYyqwd7WybIFJVYJ4FFwXzZ
J9/yIs9NiBXcFMzrRGhAnpqosgqQZay8GVA35+vIfJJCLz55c/81athWviTkJ2V+vhw3RMrjZEKV
EC4XTGIIC5GimOq/IB3BdsQIcZUiUy5RHcQAFKv/k3wp93SElogb3JzkS8Bc1yMOceN+vx0dxC65
3iKT5iSI2I5iXb/wSnqfbfflS7I1gqSJJCcSXhVFcpZUTKz9MqamTrNLWHGatlk1zZF7xl68fGO4
hmtEh1OY0zE85cPwN/S+VZF2SEwduNkNVQX9IqFsTZFlMw5K/KDzRvO8iGxXg3H6v+LH0pAToEZ8
mCP6tLZ+uSI07bANA7MUDRW0k8ZqxFVinM+RzoVu0iDCvGj851fhs2aXTk6j+pN2TsPFSexhgkD5
m+KsH340rkQR8rANOpohRJnB09WEe0ChB8ZHPAyydH93GXyBW8+7ULY9LoYwlWToM32U+W4TcULF
mgSUsg3IKHUawL5EVUjK/0SlbOkyQDtXI+uIaWoDfE9UlZh+3LN13LxIz+uLg+MMvxLTFqWutGLD
QsiJMv8c2T1j/64fkHMPwDKbkR2OAFfla0DmdgHi+p0u/tlt9OSSDJQ4WTFsXPY4mRnPfWiZgihy
0B7b/P9BONJHXWK/FXN9RHozivUx8KiA3aTACeRyrk3qisCNIX2tp7KFHEp5BmH2bXWU5foXMaGW
D33NJMiz4Y4wWwV+NnluFlD2iQXA6LzKW7TAIRXgeWGwGVmv2Z0HHoLxKXK31uGc/HE5r4yvMcRs
iNWOtbr9NAt+3uP5qACWuZM/IWEETJEkaSCQ2QCr2MP9MjD80EPwNqmcpCw0KwyFpMCprlWKypV3
fsFC6y2fqAp0KPoAFn5fsVYkrIMnRGXt/dmJmxAyvevGtr4EtEsO3ZGJBArwnWAUs85fDvVscQda
zFCBHlEAZZq6jP/1+S3WnWyi5jj8tvqo+HQEqpnMwMdj55fLPgViQcRaE1ar8FvAktzaGjcXkHSw
hmcZwNJNOGssR9rYNSnRcJGqnkIWPDPskJR2hO9hzMnf6VbHGwXjoGTBe10jiWYokoDm0bYSmOGC
Z+shU8nQeUEbhvVofaQRGD5RK53NGtb5OrRBav8zmFytlhblTPOFl90zry2C7U40ataZhlBc1n1/
wI80VQoT0DZHlwdg5ROVeAjfhmbEi2z/NZq2d/FJAXRbAreSUdmxwcKInl5dXPUlhiqYRuaZglMx
4OrvSJA0/KRVZIbjzVl++ZYqSfuV4N82GpMd4nIE6kAFjlcdcXDNfiXOXDoAJYf2Ub4d7EORHjGC
wME4zF06BnHEytER2Ps81+70JqyihNX5/p5/qFs9JJbaFK0waZj2EOw8JlNMyeFvn/PjtjxnmE2U
6olOirFpM2K9xNx0ns585zjk01RmE8gbJ0RXhK1PCPUCbFpVNgQIVQgbriIQ1LdTcZJi1TjQAKHi
ktzmanCsO8qt4lWrA/xOz9CUoJVvJwnkLkA0YBqU7gObwqKIr2hDnkemr5TA2rcd/Cy4Y3jBMTM0
omRI+n4VtK5nvgupcNYhmTmJDgyHI8c5ZT0ub5LdDVONnqOtNVuNQwJczGoVGux9qOhIXQ/IK7s/
uakAvZub76D+LGP8lSSbTPananAI6cwNRAQgpfQxFs+GSkkan4iVPP3CZgmMGLGlB0nVvuk8sWbN
ekmzzE7eDCSgdsQRa56ZCuhg20mFG+5Nd2cgzlSPL8SWQceJx5rlWSthQq3LNWMTnXy5hnRqAuMR
lIQ9a8QxsDB+kr+uF/2PErRzWzzGG/O3ZcFeJ2m8ES/LsnwHd4srImeDJnVgBEELrVy1LrnEL0UB
xxrxI6+Fn7AgYQi8S0pwFMmfeyaUsdwWlXHIOoGuFjvEEvI3yDWViFTqvrRbBhgMF4rHqL4tmGzM
pSq2cJ5UQe/25DBC5l5zfeTWkwom9O1U/ItWArHBfZkWHl/PdkyvQ6TZZLLYcJSeO/AZKXTRyMNF
tfC8+eqg8LFC6WNWcrOtMkA3zzigEQMjYXf3AdOkcgmYbKj9810+MH0WuTi0VYTfyOpZdKul28Cm
c6+agrmydJHUFgajdjEsBCTxD08E5yhjrOvgzFTmA5ca49GFxalEBzQs/ZkjXdJ273jO7+YbwjpQ
S5xIkJynk2/BcN+5SfFQBBZNx4rET/vJWirhCueY90aCvNsC+8Hn78CBonboxTyyXKFgQfVeQNzF
0vw4EfRKtWPxE4d21FRes/GSXkSpTLIqL5AaR7CxgrMBhAhn5aDRqOcCTHZ7o7xZQ+Z99rET/VfY
QTO/iTFJO1oISvqARz5F5m1vg45eBalvUoo3qYo0jpc6AKarvf/unlymvW4KaQQ87iJjRXhy3SL2
wL4pbkWrnEhjYcG3FU99X4hzyzi7ApwNguuFFvnZDKQOuzQixdWRkUEdrY4AyGbW/gU4pRvDuKEY
ouK5iFTcvoV+c0Bo+Xv5Y7hbQhsB/insh4HbYFEWzIXFyaaj1Wk4m3Wle4uLEIR8J9xmG7oCXMwz
7Dm/64yEQkb0WtimSNw5lZOddyhi//9BPdrqiZ0qIp+bQjvvidrjOXBRyZJvmElEkF4snRX1feg5
/UqauEf1PYLBeuDQApJ1jnEymFtmx7pCwsUs+lQqTNDEz5h8bj88ttVq+T8ky14RgZBfx/znTdOz
wewoW33o4LIAnsdTUCUBYHAz9JhKhTvag/aYyJ/pMrYdp+a2zSewihddFGEKPeQr/dV42a++fa0M
4U59jPl92QsiCnsnmVRQlI7E80kdvAZdoJdit7GAGnuzOUetpKtqzdnVt3Bsw8YLF72hOmxWWByp
2vyc7xNp3PfNMCunCij3zf/alZTL6FpXPa3HMvgFYlPTOozMXV8bsrGSpEB4SLXxmMM1Q6oQHi6a
9i7SUsWHChtthk2XlBS439piKssw3yU6o/MxjZJXfyd/cjOilldPoVUAG2G6rOkBf3sI7DFXZkPg
JeR5Tmc7mCD27EBfqR9PIwb/1ydr0tj1gMJ9fbTsZG8tyhJXycAntE3arJ0mmu45aQYVrHPULtBN
3jXUtinC+aCLnYU8nyCCDoUQPprXGs0+9PgtDHw+CF0Dm0fR7IPQS//iMfHBXJXskR+xAI71bZTr
jT62SscfcnSCwG223+iD9ZE/+sh33e9X7kNVfsQ53luxU8EHGrFsqcO6IqgCxl4ELsPdbkCmjogf
yazL/vCqyeDh+n2TxNlamH/f77/eU35TQls5w9T+vAsaJqtxNeLM4j+8gtGSNLbsEDRWu/xQhoP3
x4CqdP5gNPFVZWLMYktegfuSILx+81ZreLfDTNgDnPLvJshIl8L12tY2sqdYCXgLv5k0bk0fjl9f
TSnI9rvNZ0v+B7vAfvwph9OeufLD5mMDJ2pJ5qBpF7QKUKjSDxOUilQ3hzrObtW0tHqr5AAPr2Mx
H+0aosSsm28Cof2rrSM5DwolKoN+f79SmoA8CSn8WmBWgzwI9YHKgtvk+4ZwMwrsKbva7gFwjtpz
YY+Cdje3UNbVYvd7qJSnqIOSSkuxD1on2vPTXdT7/mvkVSmmQity2pAVoQhRbv9rybLik5OeQkmk
meKVFFh0uqp58mBq1jnfPnNe7tIIbIHx/VMf6QFs61canyMc9NYHfHN1eFuE8RzK3BGh7Y/R46LF
pVud2NK2XeDRdeODftN3fddNagAwSwP/UAwFAdAtgHf4UrJsB/0k0PjNKLUamzuSzhM4+426OAhO
EneX6yrKL/F+a2esyUkO6/NJGcsqeyIWqQ7YkBXyt15r4n+uPIgEqdZvFDZCRGzMo5jri0ZrjZS4
f6x7CjEqhvCU/P1iffREIG/sDxTjURVY7DKUU5wumTQwOLAgiinmSNNkpkXeYJ1AgVLlq8evg1qV
+PIlV+7Y0e0hKwWRYrvrtnzAwQh2ly8i8msuYlLRgJtBbkHvDdcskd+6ptbhQvWn9AV3yzXkt3PA
hlZ3pNNyy7xyoVuSVTn1QW83o+TkKPgrpCJ5HQzdreFVNrXdCMbUnUdT5jKAwwPlgGj3loF3Rh5p
vCxtEBO/sKziETcjCx/7ZxdhHrREPLdDxGA599Kj/higlZsheaR0JeDBVFNXbk8WKYIuiCYkxBxF
XM57V6RZrnTn9BFtYOHcjaekXS7MGtjsrYjxhTQO4rzxm5OQZAyRYU2hidJqiR1Vo9zdP5ZSIoi6
uwlw17hFa9jIFKzWdnOOi3G9TPAka9EEyJ/VPINBmlq21bDjEH0HpS+b7hkhxFz89hd7hWpGfIxg
EDPL1BbAaiMZF91x07VVl/l3ePtdburRKAnIKX1Ku1Z7a9hUcqJgLRFuYpMD/dtJwTajBAtQ3/g0
0+LtCJIT9Iq06Zx5mH1Fdm1OIhWiMbUwRlELxpCZMjfKfBcK+os0m/VqXMswJFSesZm6HRG6EI6A
1WNDociMnrShOnBffFF/KLaH3DEFg6rbAo0k4Fyr90m2rOK74wBKNyIjs8K27lEgvc/Xxn44z8jC
arOx5WohqPFMIZDXH100QBhJxRY2kxAeFvi6E2Xlm/oMVXDMJkUje6hgva3mznmYrhZFp2zKI8G2
1L4oC9HGG95Wi3h6V7BRtMQ4XyDCCGTvOmqGP2yvIXjqYkaob+rgNJ2jEVgVksuI5U3u1+avphaU
7WhNHxKEp2meZENq7QY+WAX5mqr8E7lUoD8XO0E7/sNdcuOL2EYBuy0UUQwZW8HpNQP+a7arsO2w
I/bG6wr0wm9aFYr7Q35HjFGTrwDTCicQfBXQCbo/7tuqxiMHFWhltR+xrnX4KIvT9uOYFLuzzZ6M
VYf1lPyXM0F+Uk02wBUPVQYaYw5FzrSB9xn5aGlmKRlYsk4TQv0UoW5VyoCIQalFcdr0lRMkFAYI
S29Rp6o4DPbnfotj4AUArWW7GYFamJdX2bS2kxbD7HVxFJXF74KejSGlYWdu5bC9AKZPkYRNyEsf
KiIw/u92/Vpsfhv5sygOSOqkANADAbQ6RoZovuGDnAdQV43Vv61JdZHIxYKIgPZ2hKEoBkXvf+rU
De/YjdhXZW//f4xWPhCf9yEshYX1CjxfUKRx9Yj6XefeV35hX+9Qa7TDBw63fPj4CHOunUXOm+U8
H2WpNe0u2KXQcHnG3pqEXUfglResJfpDBfQDQDsLWxZWoKdjlHgDpM9RfEf/2cQbGx55K90xOVdk
LzK2az9D3I/wHCjlZJxOzUyca1pYI9Pn78YkJYZ5lTfqBY3XSdyK2rK+0Jkr40g4oJb/LXIMj8Ua
cjMV7tcsrtJSeWApKmxawraCyzboFhaJsGDMjs03MWzn+icsMxgkndRIX8knoBAO6/ImBSsCPal4
neIG2KJzb4c4VMZVtDrfqdFspuHKE2d6ZpWiXzxpa0UyoCS04Ixl4/dJ9oH2G/QiTtZOqjxoZ8JI
ppoVHa1IcDZkxcK2q3PTWvtx0AMuB54Lqx7zv3gvykNvjvQq+/H/LqMYJglLB7x8REtYDA29+e88
rBACUrkq/hfp5oqoAUMj7LJUz8xDtgfWvSoPSBKsoNp0cXPM9RckY6cjFsuDr/T1X22Qs7gZCeoa
8gXjVlADMb82xuRm1EtvB40VmCPmbAKHK7r4lnb0oqSyuCRVEjFXnq6CuEF/V1rVPNzMRCUB1hRI
skChPQbAaupRS+wcMxbV7DRyalUG18pv0bKeeKlVBFZ9JSveEQRO2SRah1rQL6fCNRSZxTPQ12mD
Uw/gBFM0HdL9UEHxqXDCWXW5/q67J27HvHmb6hjzW89dHTaunjTOK6fSvsOszXZk5f+joWBDFW4k
fgSbBOvmBQ2DDaIGv6usp+mQl21oeAXydwUZuQRbFqkqHwFSfOkhf2eqPvDsDRHG/bQhAUcghCAa
SU16MUorfT9W1QFVRW/e3H95seNeGX6GsApau8WGLgE+E3+UwnNBgiWKYN6PijX/93xkDjxYPw83
//WAuTx78UcrrFrYFyws5Ok8MnsFofxNy1N7gmEAtAKpt5ad8c5Rai6doRVFCbU0+G6CM6H3X+aP
FFqNfsr5119n+/WaQLIIYe+0BzLFkh3WQIHOWKONNQRtYW4igux/e0QRgeqoT4bvzdjeegJAEZtE
p97nd9JAeOCC1WMIuJNhjNvlUyKTl0ZJuusBlDqVq0AF7cgkv6fm3R24QBFCVYj09WwZjhowN1Uo
6y1vw2xkRGts/MCzIuOXXcgqbDlLWvb4xNcJEURnlSrx2KahV85rjBr/vOvn1rUwx2utcXIPqv37
NBVrajdLb6V1hw869MbtAvFGnCgE5QKmgVjm3hXEIZqKHnS3+Dyns+rHe3NHRBYQQJwNGPiNGTn7
xTqiJRa2yItR+PspRvW7d88oGUqLIypqOhjY7D2TYC/tMvstV3qeDxe9ZxB5Hc3y9iaFbR5nIXbQ
KfG9MjrMZAQhkrXDHqSZQwNLYnXL8MkHuZmWLssDTGK2WJedWPcdnX2eVmhAfcqO2/FpOXEnUetb
hmndec189fzXw21DSH8L1Yb0EY3e1tbEEBIPuzkHkoqPW3/btfTgPrWv/7S4yAIjndqmL1cmprxv
Em9UvHBAghywVqrf4KuuEJIFyGJh34T/fqpFQPrXcXIFiOSQT6bkRf58VKWhcNHgHoSBeuRSf9bA
uWy1MEWA304V8SJNMDKVHihBj2LTuJS+8Jb19BaQej0sx/qgKX9LSTcf7lx5/xZca2XsO5zyekhB
r1QtWaD3DCxF80biLLB7ofRS3HZEe4hjz8mE+0sMl87QsuSAaEQyCQv3RMnBx79kYZqX6ES1bF26
nsZTtpCU/Dn2pAlzjmLZEmKLKwWgCwxxkQmwSp31VxXZ1OeJ0UeRwI/CJmnYQiqSpAq5XjxK3ILm
tghKdEpQk3n2RVBYXq/IZ3E902c9pnAYApD6B0efv6AIIBVxMy8Lfa2BnopkH11QFHF5Fkmlsdd6
Qw44btbfHNlf4ngSoY70ldM3DKRQSzhAVfJ1MGzk41WjRnPa3qL7G/+m8DDp5+jZGe6n3ub0esaj
7FNb9+R9zZmdpVDzUejgql3Hia/E346BQXBOKJIB3He3MiEFtQSJr4IdmyjzuHGHbOIPYV9T8vTY
PiFtb63ta/U1cicFEY9PX1UycXxxTu4oiLa8m8ovhyy4ZYvYuvME0rPv6HLJJQQIeYllKQNu/nRJ
ih7oYGPa/x4DKgookK1NoDP7Ep+HWbY4CuncY5GlOWKAwTaVx+W4xaxtGCFtFLttPLUvVfQ0qGXV
oMfrab6wHRkCd9ym6rBpcSZ1If0UvboOXamu5gDHLl15JL03Oya36K6u5if7wHOtcqcK+jgdq0Bi
ENKVthySNU9yB/QGy7VM88iscoeRoqpAQNaqoaVJ8uUjKPCybKaEnPD2+HSHeXyN4wy2/JUD4RC0
te9srEaOE66whCwR+ug/gCfDpUoMGb9LE5BZIbkHHfBaPQjC+ZWbYPQD1EqzxpmmCIErQJ9vYxoO
S7+hnTgv3Me/W41az7ookeFJMFDuPN+q0gLAQ35/zvSYcMdlD2x9EBEhPjZ1oM5GTPoep0Co5OCl
u/hEk0QblPWabcTedpSKUB5QlnFpO1Cg9oDoGZN8J+2U1gXFdVqZQ5ZApOPPtla3Ce5e/e8PWlDT
zNLdbL574ovrq3siH8JaH/LGL5RrhQ2dmycTTucBr6gww27JnRnsnC3mWmP559WbeDthB5xSFycX
/mhIYNuD/n6wWZb5AGkvv71b4uTEqXbw9yV2NOzEqKstjXMi/DGGG84ZA8gDdog330F+k138aOmF
f6Hkdc02+zxv2XeGPM7T4Duicz9cazZSojyhPcwl4oG7aWJBcMd50ZXiDlNPBE/L0XVptzF13cc4
NndPymeMxCp6ysU5o6Yq7Y0jd7mJ3PKDqc//p8+FB18suclVCwZGBUVsIX5UfMZ9agSz/rlRrELO
HjiPWzqSthuSs74JJigMH27QU/zb1McJdPqJHIz9xqihFgpjShto/Bqtw4zq0PJPY4b4KystVRhD
VppAkSVEZpunTZ7UAFbbwe3lFNudR0IPyTfb9fmjn4pE47cWslxkGOKuO6mMRdX8WyZSUyDPLuzI
aen8DSZGF6uOftN2+KJO7bQIn9SL+X1Ib76pb3STCbsy9vRvmzyltS3CoqifmrfSNAvqpRZT4y1P
qLKgqVp0LTuF4swmTacwNv+txHrUO7Av9CBWGWzbWHD1UdHF+mnZUK9Uayx/MKoF/e+KidZRzcwH
Btp6Lj4UQUR8Vkwx6T8VQcZV+uJPpLfefjoVPW5CBC2Tc7D7m/Qtn39DpFvHWNWAW9EhEvgj3N65
Do9Dirkol/x5LIsov7hsZYGj9ANUrzqo9/Ctc0YEIRXgTOH5HBC8NGfyVJwfCcLh9iVoVp3g8RDp
tH3JBr91klYlrg2G0PCv9JTKa7KUuIO2IAydB0mrmIBRXurj129arCAElpPVXUH8KGndcZ6jZ5o3
D3sT8qhZvRINL41MB1+9CmlJVUsKlfI05hlH0SFzVEhwdMDKCKBoFxWoEF0kVPB47P3iGsizH80W
ai8tESayOPXepLiKb3PreWTj3m+Uaxx2ygtMnLv00lmkWG22SBiDNuBjgi026lfxvtF4M3h5AkLA
We81WVWFhLPRpFvaQAOqGTJNv19ccVvfu4l1FGGgcOaQtgUhN1viuR+PGYLQPM9IRCkm8GIJ8Msv
o5uzQH6quAxHOrHWyPT0HsxYCn5lwou/O6/7zhLMkMCeMKU+HyBCpLnLMU1mTm/vBoOWOsaWz5A7
xkB9mlSCFsvXa+Plee+k57jyuzQ9rd85VkCeuU13Zk2joYsrjuXfxtWgi3OWdlGztRTMs6WnRcvH
7QHux6f62IYUrblF4WtdON+45rQN8kOtXmm9FbyekHMPK9X6D+kpQizOitKd9TEeVYGspR62WkDE
xp031sQ4KLND8L37i8Rkd4q9oZsbMGcT1gOSQT3Nms5+WRUpS1mlRlb/b6UV5JB6XFH21cOh2o5p
nOmFWPnGr6KMoZHWAWclzkAAg5j442yh+RKhQBfVMYKbhUt2AwgXjYpTB+BwHoL1CwkoQSRVBViz
qz4q2JI5sXuRGTeFyvXYeJutefBjDld13S+MJneKQ/nFis1J99W7tGknQXA2BnkH2GKlfrHgGmy7
VSLfY1RozuckaijZb+x7Mte26812RznYSUHgnlusSUJEzyRgXh43uMZ2HvAiLmhbNoKNZ0OZUAmf
6MWwtTkStToljw+Epd1QqMeaiLECRecdikX41fgXaxNLhsCULXukIWLESG2WQDu1bpk8RocyvoYD
8Crv2UCz7IOwoR8FbOPHxoTGx/Jmote/Aa4T33dwxHJ33G1sCKHxSN3ZjHgl8tjrhlJlHXAo25jg
tGWDVbAGA42cXQS/ZvCQ0ss5TDVynGyyjXDByCx8kZv0YxWtCoOt8DtqBogdz/pOc/SReScLo5K7
bcSROg4niYZWgbR2TtUF+0y2MmSQtSycwc0SVDxlTpI+0AB5UVTWnPRJnVPx8gu3mZfoR1VzPTEy
aMN0UMArJBAIGVwa4mYEcpMXpeQ5N+tY4uxRzdx3TKY0LpjX43KnkQvlGiONONWfhhZjAWv0TWNn
kic1Ap2DKNZARHP1L0SSCXKVyK3RgHYBHiQGX9lMrHZdeieVMnFAhaXxqGG4YNM2N2KQBg1/YjGS
JuK/aETmYHo0g9WuL92T0fr5SGZjM7YForHpgFmYpOS+vTzVNCt+IMQSSaOAXbcvwX70DzUDgXgM
kY98SyWkiRl1GLjyoeuQXtzJaTtMFMSKOIB7jBkPA18jucXkZ1tBSDybt3zYC49bz0HjCkPlZmqX
qeIWsq6f3TUgPP94qpIMuhWsUh254RsxdI4gWEs3GKiC8vmZkle+0eAgLt2XeKis4HB/450uuKIo
W7Iv9+AJntT5J8at1MTiO/Gif+B8qpnGoJVQC9MAJPEmjiyMuVH8/gKUGh/JIy0kdF34prQ1VG9m
TiI03atNzrWTB9h0LklrmnVTIqyfIg9U1Aif+JNEjRbl7YpdTiOlWn3UwQMl+CsEzuQBuXsh9zBj
wuvOuywOBe4b/DQeSSYxUtq0IHAS6YaZYrhL2C+0f37Gh8Mtx4qyP7088pC/rC/Oc+Hgnk0LFyAB
ggqBX1w276H7r2oDdUTUkZlsJihBlbcxMzfNfC6gvuDFpxDLnYZ8JoZ5UZ4pY4R71iYW+6gWESiG
UGzTiulICQ6CKcoZyJflRng8Nqs4pckr48fQigll3OGJL/Kn6wdRDD/uqhf1qg+efMaYjLxiagdi
nRLSjBE0K9bQ6FMdz+LfGcXQCGQyj4Pu+4YKJPwfRKGL+njc+ekT0gYL/zkIp+Za6t51wcbfiNMV
rO6p+sgIsw6FXr4vU17U3TVv8uyMjbaHZ9ns6o2jDu4PlaJQmNdbxI/ExLW/TIcbwxTzKCAVcmLS
kN5gT44TRxNY5gNR9shYuba3HcHajqK2Flp0s0vtqCzk0AP0sEyNspxDpBv/InQFHuoaPy2zS7mI
RNSztpiWvMGl26FLbLwAKgsd7TszT9NqmXmbSPDllUrDLthXi8nJ436scfAmMCpjr+QXhVndNydr
we1+uiwWxzi4REOaqNMBD14IgzKyX5OiKJpkApJeonJ+iAiLvXw+jmOLdQnfLjYGLG3H5ao8BmqV
138mDPxVn5oOHCRm6V61zAVKN4/XKlUDCMkrJ8CoRZzmaW9kME5maoqohxRlAxTqBqZGOPuTkW7o
c5y/AYnTZAQBNpTzzGeYskNDhMl6X/BAAY7uSruWfv85EBzYA4NFrg0pQvuyHE5LiyAAPLeMNqTN
1zD9y3a7lqFaQIvEW6fy7wkQ5e3XD/dLiU76meNwDxCbuOSE1to7E7Q7HbaWqANemz+P80fN3KjJ
yjY4roOScNcN7JWx+2eOb0YEBuaN9NN4NAN41nnfhc9BaUdErGHeM1PxqqvvW2hHyIz24dO2wQy7
pkFG6zlhPmWNlPOf6Gan1GUS2E5QJJ11vMx3Xc5yfiQFdghFhiFhimxsgI1aKRiTxz4gHUvVKWKz
PX1b+x7HN6grf5LpN0q8NcBrqJU1j2rKOb/6minasCFRzsaPgfkEWD+1M9YS6ZPvGEoyAdgC+mef
DOryfb8sHSVNAcjWFRnmd+LIOtarHw8yQeaY/TpjLPBPjhkkCxl7SYWQ2kUo3L4LT97WquP1+9TR
4bH1UJBcac3MWInu/OMUyY8u+gBNN9diCV4PNglDveyiJ/8NN/PUmlRh45YJ/5Dj3kppMEin6MeN
O7rMWeSpMMGBSSNULi4CC0dU+c8IUSdTHY8JPXXfeI1wMkYxHlKymY7Q3GIT9JmS/SO5ReCBezou
ZSQ31PThsVicY2p7uxe2yzGBEvHT8RsA7jeVjGImIb3QWpneI0qTCJneaYNLZf2AoTVceoZSr5nE
/gITAAbMTLI/TWgvAiI3Fsnozz2eegqakWRLF1Z5lh47JS2RNTFmBShJkMIOdaECa4B2LOvOifHU
7vcgrkgWbTpXp4PgRkzdbSq/VtvOabobd+ChlBd3i1pzdaWN3+jZNTN/i2LTBSxXMuVJ8Ky4ACYE
JJhEk+cxdh3I55GbFIXaSKXReAJn4OXX7iFn3G88W9Yr+cTycdDDZ6BCXVN9je92QqEwXETNf2NV
hCwE1HrkRYrKwPXOVDi5dLG7xoJg+hHj+B6Q72UyuLgBGpZe7idOTwHP6HqQyPteL7+5BzDpqe0p
D+sfoyZ/WCx7wvfDqB2oX/rTDJWpuqzcgaCy+rOgQN3MvHqBrGKgRQ7aBSArB0JBF8G5cqSMWVo/
guICQ3P4YaYRuruWfk4677lsktlZ3IUpNDVhdp/M8D4G5S6d/0EMgdW+0xbndqfQKTV0QTHWUW/v
FSXZUGcVqQpfW7M6Mje7nJzpJRxtfKMHnq5qyX6lwJiWk2ZUurJYkstewzwHkSVg+Cw0JlFu+vhc
toTEM7TYYZHOdV426vhcSj24+IdMhhPAccQwNMFqJm/qmGdcjN8BFkninoxB5wwB6kJzcAxxS4tk
7ldRCGtsJrH2fqXT0Mkrgd8fRNbfLAw7tGg9AbaUqJFjfvCXk1uJ3bHRXnJDp/c+kYuMGTr6YGro
v4Gg6VGG127b8b9kiUnGj1XipFI8ag1QCbMmr8Tny6NougdsZtSArMOhaTF6NSSLF5hfgyg1Asau
65tL2QOAsBtxPKy3TXaB6mILFA8FnIE6fdFpSS1Tgu3OLuSW/10kv+ZAoGrOllx5170Pqo2i0QIf
q0U5QL2ZjbP1KC7ahgzl7wnfPWSeO3I9K41eiMu6CO3v/Tc5/6xTesqnPdWlm+WuUm4jZ2Rjjs4Q
8lVxrAReYDTOrWu3v0hyc8+5NUDJ/F3tnetTUQpbZPP6TeiDaGTGuWDbHW3YXscb0GfVRbeAWKjo
AFFKIKLcBoBWX/IN1evV0NlqxxucQknHDC6++kPlTzGi44K1NcIvAMNe15esdMqiObhJ/vSYTKEy
cp45bK1btuX7kPU2YcaCgxx0cCWI/RdAwQ1Fo6Kl4x1Qc1KLAr1mrINDmQW2/21w9T6oy8FccMlx
hZAH3abg1uv4f92N5oU6LEc+5w8xoQRvtyNCB6yUGhpOEnHAasyC++dL8yTJ5UNg4JHH1IyLcbie
Dqed9Cemi1fm5jJqL/MSjKS5/bfBbHYzizy3YHXt6R1w+CkYlpBOBb89Fdohju8MTCgM5wv4mrAz
MoKIxgQ/NRJhGgVKfMAj8HJ1D1Z7m3xDnfTOP2+uuwObMVdSTFif24W1hHUuGAmIFL2YwoRiDjiU
br+NJlGvUBKy3ygGbvMGweDw2IlOFL4jcAqjuJ9sIr1HzduaXyHQubJUR6epB39hSYf/G+70F8s9
GNY3YJQjZQhjCYGHl9Stao1j2rdgFQZrwY2Hnp5qEgNizd43eD2vB5kUiVNeGU+rS8LZwW5szcXB
2768kt/MvK6eV0cCOLwFtfNM2qwLg+0o83xCvMBdN6HVCsNe6JJp6ziaarksFqduyo3HjQQZ2IuO
SyegLu1oxxULQl01ghytC0dwG0csGQqmTX+XsnTQP3P46oz8aIxgXGifa0Dw3X4k5fVwqN4c8Qu1
FrCai93Za/4bhSZKjQ30NuMa9QmEyX8jahdQPsWgMibUYPr+S8D/4xxdjMqpZLE1IGrDvB0/Gmby
Tg8RCmlC54yWlv6zhJnbQRVe9oAyVM9YEnNJV18+Ves3g8/t4Qzqf/jQlaHzVnFZMZXKX10esThP
mxDq9t7ErD+ri1Y9NwQa7TwUgkfoyAZbxygVgb1ztpOldisKOaQ+3Uq7Zep/rkM4qc/iUYmiv6YP
vg0+1HD36pnV/j75atQqwJE4fPWd63O0xhn/mNxpyAcDg2/h1GHx+5HXqackmQPpEBdKtnYzHj69
yOAAyWROjpi/jhcx6k6fGp3zYCfbdFXSigls/sTJJV1EgW6Ux9EhBlSbDOcu3v59cmtzMk8e4Uyu
BbJQGhvv648K4MB8HULsFsm3y6kd6+5m6NQArBMwCATPfTNefD4eWKZKn4Spdfh/qbLcW6OtlDVx
1pqCR1vtZt+uqXG9i23slOwUg7W8EbhVCp71PaIxgSeVBoCyj8NYPEwqNSVOd3P4hcN03K6xSO1r
LoQ94vQxbuVehvpuuV7D8NhKpU17S9s0kQgAuyFXoEWzytNUFdVzdmg1nh1PSfYYsYxkLZyejrBF
MX91E08mK+L8TK44qRy6ll19DCySstPF9MgmA5a0F08f1SLoS3DxunUwVJWf1eeBYDJRBE2DP3Gk
7H7DJXatm4gdYOct5KiuBw6oAX19F9t2CAKZ6Fjv/wzUFmS1esAWWWRONLQCdkQiUVp05qa0J6Fj
amqduzBqw6vKxItWrSLOWA8uXrN/YINuRV9pDjfBB2r4oiPbXuh3PfdbdUDxhrPiJZNQQukc0ozP
AdACQwbzIg/CMTmB+V81APmq8ml8iYBxb2JqMqzdNhCbEU2ic+kEE7RL0Ev2zkRCJ3Ok4X3iOGcP
Vl19+DErtXuqoFbHiG9yjl4EsaZY5ujUqLOslXJdy+CEHxC+VcV4Zn60MI0oH9sDynh/+xMNbbHK
sIcwCCk0dkPG1Ib2lxppIniY3DbsCHGzmnqtoxB2b6usPWPN/Eu7nFrvKSsaMh8AWXmzW6Szm0bo
wrBDjwT/9XLGc2MsfVOPFiHTkgBBH3Zvtn9rYoNrfB57YO2+DNdVuLKOdl0gDGHXBd6cQ+LJk0RV
YjhnnS0JwVXHT9WbMqYvcuJ4KYpOkVDpAZB3Z4fDp3Zwb1t9PJDrV5Bmh2LKN1Xu3GLDt75btfQ/
p9uMiTAc/KqQ2KxydGMhh4kboRihJoH4cfyBpIjiFIo2AWHk6Ps62DMgYgvfavsLvPzB26fX0yWp
jZynpQmSjPicIqTAfjgPm20s5UeEHAUQTRYKaTLctTCG7GGmFuq5DmcbW+pTcCJLlrn+tkMFr/Y5
pqdMAg4s2HapVSE/SD/K1qmAXvJbXH7ILovt4uZRzCSTZ0IKX+c/vxZUleevLFGFghhqpl95HmNE
xHIXQAc0dTMgGL4JDLK9dgduiEGfhY9Lr6aJWLsXJEMR7JZDaiztDJZHunM/yfXlcEEIBf5o4d4v
CVs3mceXQ6HNE+2rP751nQeR3AH2Eoa3GxC6UQeZTckAmkQKMOsACBTv3pe0wMkp84TKZsjoyJC6
5WWiBR1/KiZHdGyeTunTcfSK6rjK0XcqejbqIJnyJNntXMz+ZIHe+esTubMnKM8QdKFx6+T0fo8q
NxRrPWAo2fyKw2voIvaeRQCzSYNKwEnyG7OrwmBCGOvFGmB9M5ZcjJyIqleo9eb+RuF4byPTtR/E
uAkj8NryomdCSxqY06WgZfFDHjg4AYMNjcAalyAnHylFWQ8QKLZu9yx507ZnIJPH7rvh26shwJvV
IkUXgQY88kemZpNJO6FIFiDlZGkMmaUr3yMQWoke3bs8WO97ke+yi9V/XvFw4SEgKOwHKTBfKFvp
zzzK3KQ8uiBvqUkdQFZh7lAWHaslG6PiDvm3tDbzCyFPA2umLQ29SjLSjVSnEzn5EDZIRSB+RYB0
YNCqFM0yBFH8AmDbMrjcbadmZm1QQlD1GzmcESi0A/C2NOrRD4sdgz1+7j8JyVUj8YVItw5boeaT
pZohhyQ5qdVgPssAa/XOrfTolNGEtEGzu4a9cnwCtsIWEfCCaj05PkXG2L8p6ns96fePlxMx7xXu
Wyas4K3MVJbnyKu0iAplKL0n5b32iEPH1I5wNezNAMP3DswXEQPojxb4tPhzpq/yBVWlqtWjP9bC
4YA7E47I4VAVznGLpSL4CQ+cbyKIcvJEpbGmDtsjPKCVC9wJH6BWDWZHwMMZ6gZhaHPSbfwJxkax
t9DDqa1vTFNbUAH9E8CZZERSkceBjISJ0pKRWeymuzu4I1AtU+rPwAKYkI1OIOIo7Q5lWBr8g6BK
tUatZ2nj7jnFeHEmW6mElQr+JqR1lpyql/3E/97MQW++JANDA9QhxotLrTVdWclkWMOU8vgZ+2Em
uSqEyYyE8n+VX53C0nDklJ5O1Yv0iW5n9MHJk44+RmP5pZ6qAeVryBhOpWZvn6TL8DsWsUHARXfQ
cyInsZwH8FSFpAJ9jjpddgRcDrJFCmqgYjYgaqZPpgDBz/MlhGYkD/N9GOki1tf1Rc4P0Ft6lC34
eRLDLoeHUbDCdl4xVb9EvcNM4GGWk1KwnGrgbx0WlJ6SYlP5P2bJhUOmNv2wtcKstQjia9Sv1+dc
yk7HeVrpoT7EcOI+9jLNIOvewuf1tAQcB05YzjWo1QnONM62hTCyDCtRqQj5mlSUONyNhxNmCnpB
I7iY0nftmyarq75JZ7phU3PgzJgSnvUVyFuS15E7RXbV1bcsKd+R3GcgU52yuVJRQ4gQlhao04Aj
QePj6QRrnoIYKr5SEeQZaAHO4fMI+Bwp1GbMxYMOQG0uhZDygMWDTZb4Y4TWiYjE9ZbPca9l8nvc
/YlgNocKgBtI/Dw/L/+zRFCITA0q6Dlg+N8uc/wpFpWe2oNt0PnjxsCtwO1rTktjyEX+eGrylkw2
yLsB0hdAeiDMM6IZm3fpXqhTWvleXO4IzmgJ/IxiigcThCVgI+Uoi1FRI3RVL+2W94OlKUBCAnb7
khlZIslmmlr5kNskQkZB4SL+EiANkQH8Dkz+9kx/GrIGb5CFb0xSQBvnc86XTk4Z5vvgnv5vU+oE
B4iZX+a2qy/fodihDQLZ9C9UJbpzT2rIlyzFWPtGaybjyG4AF9mprqrRiImiUWY9vON/AjWru+31
ct4G1g5oZ3lM1/yzPYbU8J5ljgFXn/ZbYryfX/7OLrjR1Pu1LGyirznH2drfvxIMB/kC+slbywVd
aWYVYPBlExd0Fkjum+9nlCByne3+EU1cX2SzVTPKJAmoewtGd7UHihMyaOYstX64cFApYTJFS/7X
xzVymUwsbKCFm3lfNtCXqlylip7CwLAuWMIiQozEXM0RiJC/INFcaBUpHCy7axI9J/PWUjc9ofCM
yAS7i5sT9dSFsgqt6RMUgf311xgHOm8pckvBdApcBvyWaId/zgCgmnropdBWr7LtYHOYvDierwm6
PC/87z0VQFGnvqIO4g53ctnfRsV+lkjNWDzdlDbPC5GbJmYomWf7NTAlZLkbMiOG693hfKb5+GIn
xLyBqeEFRtPnQyGRGIarWFbfH/eqV2zkxb+iRxO8V0iGQTQUkGh4T0zTZmptsPPsqCLE8wJBYYKd
eA/tYHGhpcIzu9iVwHgvSfFEkI5mkEHlRXPO7LcxmYDhcHv2rNx3DdpqyQkYg5YO1YD46N2n/OAR
nJ3AAfkaHqy8hYALzxKtFyNaE1DEC+qEc5EVgimdxjlnF08vTPsjXYfzBLzmNdQJk8VUY34jRO3X
wqahMqybEFbu24U8wTKPH9h3A6r7sgDiNbVcxcqJE2IJT6g57y5Uc5pvek/H2APxiGAaxPf7WzMV
YFtN1zIj1IfWRT/vftiLm40oCvsreX/b613MimsflT31gX1zcwgECk4A6EMNkUhj0/ils8TM4pha
P325frmWUaD/7kyIzd7JoCjmwQuxZch9/DX550tnHeBIuIItDjpg5k5RWzuqsixAPmRYG0R4MH+B
j2Ww/Wb0tIQGIoxG+LXAF5gmOUFLXnqcSHdI0QSoocSAKPnZixaSlJSMpI4cf5NIhzqmwOREPxdM
SN/LrYnV24O+dKwyRi2bAHVHR/2S2bDCt1XBmY9vqeuZDw5ppVS3c0+MTiKkYCEGd8xAXN4Ttoui
ZQX8lPAopDgEFCAzkQvHj63YzifUP7ohMCbxg7DDbRynUf3pilpzCe6PlH+Cznzy6dTatwUwnbpM
DU7rCqbCOqxJwX3knn1pX4M/v+n2Ytzgo4UKdS1m8oLiG3tehJ481ZffhpnVWxKXHhBuQhkuT+Ah
9BMF3iCgMuNaA788PeWfOl/DzyewATYCgzvRXfFNw1VN21YI6qau2mlRCM8w0V6V/Tl3CPHI26Q+
3YAzcaaFVBtJv9/mBZG6L/SxPmU9/1x0HDU5N4x4gsxZ+Uh2nvpwrdcBJycZM5FqhA4faMoj457V
1mtocm3x2PjH/sRjuP/YRutI2nAF/h54V0z8QPu1y/bGeKq4VYdkgEM0984DUInoU5ELWVtrhf7v
cBWuUwm7N7mvEMroh6mhxDr85Z2wqEFn3DD3ZLRtuEi6OuJ1KOyQw+jMNolrQZb0/y5xwEOX9YtV
01OwzOjQe2pyAzzckqF22/Wyb10KcLb72kFXuoBiuEFszz6e5tR7L2CaTVnGSjleXn6Hc7CAVOhj
Gk1Hb+p2a0xlz8C5m8G5rWbWBZw4sNkPkbAoPZ83yC+m6nPe4yBIXETPhblU44JDm/fSXHKbR5RE
K2t+tUXnB2y23PHX3Ln/2TaWYj6K+s7HLJqxiib6JHK9AIqRuapPeTE6Mpo0bQtfs1hjQAVd7+J6
vwP0nFWwKZ2c9PHY9NverivbXT3teHbr1GjB9Da7ivIQgrmfRoDIyuEVJs6QW15wLhg0z57PTJye
j/1O7DViWviZUMrcWV1M/O1OvodFsQ3twiZ2Zy4o78dAbJU26Hzx9zeV6jXPaacOHhzUdDBaZ7n2
K4FVus5zRs7Lpoe6EsFlYxWeaPKAAO7ZBqaz2YY/zMV/KcDDQDttnSR6StBg/Othj1vzmiAkwbgj
1c7gMf6M4ZoudF1S81VAdqo4s2H14Bv9GilbgZ7uUL3E6D39Ga9BVlzjAJyv5CMwy/YUMsITzmXl
wpgawADv5iF0u/vDAE8XK1qUcw+0sp4FdD4PD6hGodUCLIsLO3e19ieNiMyBpb9A3tsW3OtM9XTy
t1eMOfJC05dfdnAL7RTJrzHQEwngohHNs1lCgNq0s2k0o7nSE93RXxBGsW2wJda2JiJa6pYFj3kt
C5EgvmHMPM8h+fkvE4dpLX1fJpf1x4i50t75+H/QsIL4VArcsoUThWejM7IihG0mzkWn+8QBNHOh
5/dcPHpLivNas1AF0w1lJ8OZf7lqL8zS5HXvfF+9QwnlfzjDrFptfn7WQWtnEdO9Ad3Dq+fa7U8f
Skno4iJHKMjlBkBywe/6hfE3tB9zPSIhyqFf8c8KEeWiM0TH0/nPuMwJ2icQ6RNci9E1/DEi25m8
K0kmGk464WUKvTn3XLwLGaNsi7cUdepFboCuRJ5fKsYZ/NNYsNA3sC36dYIUrXmCwKAs7609gAD8
nCaxOa14G4wc/1IiqKJPBI82GJ+Rt2cYry4QXKy4P7TuWJCHicZDDlTfikNYUa1dDYBK/0vcJg2/
cEdY6CxzmCen0ROk3eBfzjQietH30ifEoqYxOpDhVbQGxRslAX6DL4yKcEXIy6VL5ys/xh89PSff
2OygYpVNfySU4u5uuAXJh/rHUqKADsp+b7mlUslHWlxafpAyA4ujsn8f5EXjcwG/ySAauDkWwilB
iVLlrlIjZBBp1uwd98IxbEKaa9NF08gMNItea2Nd+viy8/JwJokXkwxGgdNEfFsyM4f+FJF+tnGO
zQLnIoIVoPYneA6oLbjwiEaTcR7RJJRR9mn4EagdYtXckbb17aABiX2NpNniOAy7wM6KpzIti/qd
BDBuI2del6rZ5FUqSXhBWQvO7FmNOaVJE0w5sMKH0Jx3BXzBN7xnk6KeJ9h11gRATFtZGbB3GCEv
+gjE8g5u+tqVArml3f0wvv6qI2hwsuSXPGhMXD3lXi3tZ2fB+AvcHrEsAWlJBOgRCdtR3U3b5q6A
Uv83rB90bOfIxu3dtHJ+xRRHgDFL0nExng1nAZFpUKNEtSmAe+NsdTPM0NdVHOEaAX0L/FSVcXJ6
+pJysum3f0rPVcz1Pvk7md+7wT4QnCix8qKF9Tk2NGp/PlzK/froN7HS3b28ifOWknjQM5Sx0lZv
ha55iTimussuQu80KyucEVPXWAhawUj0gneL7Y4UjkPNiMEn+dOWP7cgsRHKgkRG8FABz/9Vj0Mj
TVNjBLD6tnERcKTQDTg/ZmSJt3WovFhq4LBeqDkxvnlQg2RbTw2nCvltQ0VCuC+DU/r/FKnw7LBU
TqsqtAxe6tnLd1ZhqHxOmXSiImZwpn9fv1QPZVDdLBwbBpDL2ng5lu2XacEQ44e0An8knEk14cXa
bkOc9rBlgBs2vGzXGZKWfehV1D8ft8ZlKEcfW44XWvD3wgs6ENOf6KQ5zQP3O4zrnzdMdssQ38RT
T8BNd2AYQyyQgrx9T53b0yJ3fIAuN1a/knA+klJdwF6KagFC1aXZXtCMBwFOxRv43BQhNRDLtTwx
daqB1hsz/uVPz76GckDVgkm3958oJTPn2l8LjOSV4HSZ1k2bFqn5j5u2qRLKgHQiebUtvyvx5I6m
LMjmSrYjMxFTEhC8I0PPLlpsGjFpi+iqGWHc0V7PKCogfwsc5ObRkwQvm2HL2U+ONiPoV+unTaIf
bojrwGJhyLvQ7hENAFipvRIIcthEbw76tLaufMqRu8m1MvUeAHhpxxA8QptnU3QJxuXVsMYvao9C
o5UabcWE1oy/f4mUAGJVsJsRVIAeG3mN8u4sBHk93/V4+00q8DYezVN73lY+VcQHFzcdNmtvtSz9
joBdtJ5R3HI7ydyEWi5uafGEbbfHkgLDlgw1GksKko4V7gialdbE5DrZMaKcmEEXHMPryz2GNN7Y
wm+iV1fj2/5SnxdwaE+66MSPNZw46Ga9KCfLcoZ+PwUJyaaZm34//Pc0IXEYx3gZGgLShDlPR+j+
6VG44WyCAmNpJ1LaGqMdCGhBkVl8f1qsy8mCgY2uc7cbiTvKZBsUMiC32gevJY1sd+BSv7eSjBIg
tts935OyXfJ1kkKvq5NI+Uw4MIQb5BXXVlaM3LvjBPDK9Mac4dMzvOosZZYDOz41H0jLYg0Lh6B9
OvDEYF1e7IwzDHVw+2WpQTYlreFbsyvb4/qh/C/xmJfTFHwY20jXjimifsZ1oqn0edHOv/0bX1PX
3m6WNIt/pHiwo6XSZgxbbGAgJnwRy/3ZCnKwc5LCumxVZ+YY7eGQCIL+3HgwhZq23Ha9uOu1c1vO
kGPkCl9R9uYqFTIiSfroN3d52HIM6NcJpZcWALYPMdVPnq/Gguuj9GNAvAaJRTnGzkChjhHhKeQP
SM+X3U/v989WXvHMJPu2oPkT+TE3NZc3440AVQV51ezeAdxG7OFJfSZp7jgJgIkUTmQ6i8oDMMyT
xeRA+srnPLKaG6m/shtIq6Y9uKt+4RBQT1j8ZjB4aAg/K2SWWnJl1s5o+JjL2NoEaNMlpG2Bvjpj
0rB4EM8OxxJ+IVJ7L7KDMi7ssb3BQvyMN5DrgEEDNfZ2oE7ACBJgwBZwK9OPsCQa7dGTzbBDceSk
dJPdG+TcMex5EXtAmHtqIqa+JI7/KhdqMjPx0RBAf7Ju8f/qvo6Z51eHA7qcaYZuEHJEPYfi5Y37
78WmvhWobOrEnBBRfJSpTEHCvn6M44/woa/n8dlN0BqsnsyddUszonNPx0TPy8IEm6K6VkF1fCKK
Bo93+sUilbY+VtBVUkqmCpL77ZdLfAbz0wqal/d9RXtFKXXe4cQy2wzxXxMEkF1h8BfIKXd7rAXt
eMaaVZn0ekFiyCYAD8MavBfpMKsaNBhZbseULhO4t+r7y+gD7U5xUJpfKVeNAvniu3UeXZGclOIC
JOs0ZASYbF7CwE6exPKLLChsum28n6ouD3xB7UvLSDkwVYuy1MTKvii7ooBog+UgmsBkOlBDi071
qzrrldHxTqvAPKxohOeGm/6EBHv/9GKl8DIdGFcAuMRHq3IBnAAAtNFvO7jfJ7TxYys3+A1YFtEa
tNlZglMRtOwBjnb6vqxyujTfsM3AWGPoERVoWjQu3rDCfMeEXb9XUV/KH+4baD56oXqWU+2opYuV
YpJoWWUQtyuQrdAKCQaV2AlG+fzi11hFCRo+7uMj+jFarle4C4l1B7cgE4Ze2zgf2LCYcF6bI1Fz
UYbaqOpGeW1K7iR6RUYnnuFlPn5U9MkUPjafWuxYeGSlscLtLJytj2tyiXXLUh33dEfpavXecyyu
tbGceGi0MPvknSqhqtK64Kq2w7ZuL2/eg74RvD7r3vWRJ26SdEKn18tfPL2pYldmU5RAZJiwX3J5
3zYJYnjqTJZ170xz1CoElf5dQ1oGT2+j/GbVNAWoOzxBq15HAcQO0IRw18gWU9LoKkABdDgndRRX
NJ8jjLay7EDRAyWHDJ4YHbfbWXS3nrwNjVb9eyuhk9OJwjoyR47rBtMpQtonSGo2XC6w5R23Bro+
QhRvrGqAVq9kuFT2ANDIBLfc4g1bP8+b1Sssq/xcXHzPTz6bHJ7SZrLIVcCmJ8vcoOtkbkZQkGCy
we0fuzjfBoq3oj/eBPfZJ0FfKV/N8FsGYVBrb5SvdDqK1Epgr2Bj36Vlwz+DxJN0gHzq3z2XeFW3
XqfEmowOZPIBqj/UD2t+CKWqIUiu7jAp1teHzt2Wj2Zf9fAN2yDNTlSS99vya5DexjlMisKdiFtl
5QL3dMWn50mS2AVapUSrrq6VxxOGCUzdpL6AjoIvGHC1hvnXywuE4nv8FaaVilfsXW2RW4i1Koxl
ByV1d5Lrx3M/cXbb0WSe3SoMnEZ63BTvQSh8iFr2U4yIxdjh0c9caipCn9rVKnbRL6ox55WLJpeQ
KuXNHyij1rs8fwMdPAEbKHdkga3u8io/W7rVhgfeVDw6l+rCzSGxGjgYfDY+6HwE6FNGdgEoa2JS
4S+mn9HEpEzDTLyv+lbtcZXO8Zxi0ONmdfkkXxuJ5y4I2AVINKFZ7/il9HGLkB/HwmCSFToU+2dW
pgm6+kZVs5MF5oNNOBHaSNSH7V7ybYf6BRf76BcLstyEjqlUvDLWO+Sc6ARtyrn2TmxeKaK0jVcv
IEfIB36Fy+uunlpdDeW9gMLb5RI49mEAwfnnQhZ6XJq6F3yQwki2s5jyG8vpfsch8JaFuLevL2ll
X5giDPvgjD3Z3/flB2eNgSrx0nvSDwNwMukmAd4+RU1ZFTInHEOddCSzpTCJzorzk+s7c8BFK/00
Y7dv5pDUbueE8a8kWtNEkAnWHD0j6/mGM5D0oTHHIVJRS17CENYQ4QUu8brnmcoD1tH1cSfzHwuJ
y0EyTNbtbBUazGSblBPtzLchc47XtfzevvEVItUrmkjBbW30s0VRwdaTZWW8a8XsUxT5956mXPE0
j+p0FFWOLFUh2QwUdKSMfJj7nDUfTQTtBkirIWTLHpD3ndVPvqMCEwra2ePL/FhDUgZ5BnnP11td
4Orajl3kubMk7iAHMEm2SagiV0nil9WV7BkAfRZidvzOAfoU1Ugy+YmcYWMmeipDftyVD8H0cI3y
RXB9PGBHKdFq1CnkR5KvVWmzpfmJ4oGwJguOLeQCPt0mA/pnNQEAQoPNdCP8rL99hb0Z0vRbLjom
24J0P0t3W+1qXPb6KfJB+EjazT0QstcjaPybowtiqjazP8/EVlbTsyamuu7CHCTZW/At7FY5fvI8
vvj7hGM9+QudyvGDnOmOtnFWihLt9eyEgtd9PBFxgFDBazC2n8m4X/x40DR6JDI19xBaNHxj5sTL
cQdn4x3a5WOs6yL1sBjMADmuF1Ub2OadMqV36YOHv60Q0+ijCwjJbVU/IQwMTvffKBVD+bJb7/rn
9R5F9dZwzm71MQnfV1GH2XGXV+yibD7WjFvROGX1MQ+FaDxfoTQlWGGXVi0bCC9wHEBBFiYa5rf+
9/76ZGXchluxvWsppOfHgHjlP5b6N5g7gd7bbODN/8+CiBNvcoF8wcNUOt3u8e42xITMY3s2KRQM
t9k1j43dtUFjjMwFOxOxpCg1xFaLe635j3S+p1ie9tx8dbOe/7jvQqyXAStBFG21Y6X18tpi+4Ed
Q8ckfOGsh1JlAQNQT7NoHwyFe1JKE00L/5pMC7f4kVcpo4iEg/b07wqOFM+L1mLIMazmofYWstVx
dwmcrRi1UbHbXRTeGZ8K1+OCMlZa2tYQSQQz/VxMQv568ZylkZ/1QHgyOB61EsQGewVzClKFVOoh
pKUXlF/9B0Alo1tkwf9ORsBxEYRJxRnoVhRMxewba6+s5m7VdUvdm4DvSFU4ng74DjCbumPuwa9N
/LkYUzFk89GveIz7G3S4H3NPBtLRJLDA5npXYPNFfhro5tcJuYjLXHFxLNnrS5kXwKMw+QTOqBCI
VV7QPFh96rqSer8xdfy62KGfZKFgD4MS7IxswInfWOfuL6oJymHW3DYbZJ/v523c15FMd//SUAIf
fWKc0dOV4Kax4trrNiJ3meulJd9vy5nzpnPmuUsNCUfe3nokBuEasbrbnl71x8Td/cdaSigCoQM2
WJ70xfInl2Vsir88X8zHhuFTTcPSbhGKiQeY9izISAQAtCYQyeHmH1pO/yQC/3YnLGkeg154Z/3g
r6u2AeZ9z564eXWGsMhdR4Uo4hQRBP7QEeUTOnlS64/vts+GE4lkmXSLJ+nFg94v1BbopE/L21YH
wltF6XoE9OuP2Pr/tWqMPKtciFK3Fzd4YGE9L+Mn4kjsPVfdlRox/n0ePZyKheJK2kjg65uL0/tQ
t1/v7TZymz/9G8wfNsmyYPjKEAcbZm4l93ST/oKcfLdrfsjN8f9eSMVSchlXzyj3l8gz12sei4jg
HmEUQzzvENL6JzN+OLL3rlNgCFwGNr5iUcnxELl0iEqxTn4BqZGfEcE2c/zkDxqMfp1kfJZOE66P
NJwkZGNpQ4/W95IlVo7NObq5+xMBky0U3lI/doHCQ0Xx1auqLccchrirKs017pcaalAyS7pxWO+C
+0zdmMWYnrgEUxlNNz9EVoy0CsARu7YlzO8plFgfQkbwgsw8rf7hWsaKsfzjeFIA2otVaHGoOb8M
dmWqHcfR15xf+5tgpB8eS/n6kXQDZ9VBksmeJOwbHZCilA2+24K/XZJc12L/9p3G+vtnmO/Ujkjl
1SJovur+gC1a8tk5Iw74YVk5at+4LgHIlgav/IaLDa6hR3Z0O77gDqk2uONTqEHwNH30DPvtZyOb
JYdrZZVn5GkMxH3C01QObLjVgC7M7Fcz+HBynXESlrdnPnDBwZ9oAOBWNwXLE/FLdAUsOZ6foRzH
lgGXU5/Qnpk3tYIXX/UH9qyA8j6ZoEvImLkse1hHjwW3INWI7kRmaQ241KKW7zhiNcxI9EWO+s2a
nQCbaq3VqYbszgUbea/d43C2c0z34dn0CRCwjTZInoJFwFNBEfmXWojfSvBqGTkRHRRBgt9KlT7R
p2lBF5U1B1lee3k/CV69zoav14RGUvyFmmoqFwB/5VGvoP2Nw/ylLsGileHCWB6PWx/UPrh3XxlG
SA1zx5XV6xhqCjO0/4JTh4YitxGgENy6iEVSnf2T67aK6pdH5Xs6bxJpGNHQ4wSspO6tSNrl1fF+
l/srbZugteXnvxOYCfwNrjGAB8eu2JcWZVKXoAhe5/gBOuausYFRZKHcQtyFc9vez4NGUxzlBkqj
fx/A2vHF0kqfRs4w67iAW022qDJkSaKHH8/K+Z8VLUA2fnJB1n1kXVGVdMel30s6hrhLKSyHhp3y
v/03F7O7EeMHRcgpq/AkgqqaolYySsGzFtISqViH4oHtwaDr3xpdaC0G+aBwoheexo+azecDNXrd
mB8sBYb0sv2hlzYsjRTKdCTSbpFG9Ua+4sHckU1dWYatSKDutV5ZB8LfCtbozo3SgigRIIBSbroM
MLxm0HHUOjDCBWgldBBqaDgtBG4QhW9l8QSK+htwcHfDOK2/hSxUZ9AdiUzSDk8TX0qEFw3TeyzO
anBkOFyaBNxriIB628YKyIs0QryVqubxVpcq5EWkhNPTOqMIxbopBq1iyVqWfb/qaDU/PbmQB8bg
iJafANAONmLQZCzjZDQGKbSE6LSJTeuOYChRNKxgmk68tHqQQDAuYgPxSZtmC4A0xkxF5RtWqzmm
p668DYV+dQ77GBBfWXLPO3zXeYxJIOcIoBEUF6lFKytgA7/wL6E2v1N5oC/g71gu7By8UaJQAFEc
+oSnV2e1pqEtwNCEoFtRiPTidcgdySzQcLeIY40NgnpPV0oZ0SFSfT3uZlUVYn172JWRGi23oF8z
Jx56JDd0xLYlTriJBOiCJ+5tbUKP5Ycbt1QQXtX9aV0W7jzya66AI0Y2ryVf+wB4feWbGEvJtC4+
2n5Tl6RQM1uIokSIwc770+ulh/bN4w7LCq8FD/JBPFhS2L0YUfPZH82zRjVKO9I481QwB17oWLKu
YNfW8/t7PwlTGJ7+nsA3IOcKUNcvDFyfIPr7QLTF7tI8PRN4/kDoQRS2WlY83qfefI7MAOTuaULs
hHEtDuu7m+YV7uwsNm5zdI2jLgRYf+oIGx6XcKgOq6/4oNa+ggmy01PQuIc3ecFnDvPSH8f+LAtE
QqfMuoP9TKfeR0lC/912FKqGtW3/ZU4ciBGKx0PLtyxJdxWrFZ3k6OqMrtaUo0862ytipuh+OW7M
vS+ilpRxc+cstWgXC5vnmz+xT92NnPRVJa+T+XXpEQbEE+eijwqwyl2NZ2fgwjvTRUi+aJNMqpVS
igpytFfl22j+fCCL4I8R79X+VLF+ABXbOYhbvG4v33I/LSNFWBPsfXM6J8caHQthNMgmeN9JsLBp
t7pkLSJ0iqgY/NLt5gsyxsQDiGjEJySE3tNoIWsl3Gevmt3lVSgueEiq0NkgkaxzFVFfJTL/aRx9
rLxx3nmv0DGE3OTQh8rUIwvAkxIsm/ZKO+bFspxJiWEA37EF9RW8elEswgn9zfRK+shGZfJAeVAf
38/e4HR5na4lDfd88XCdue/ye8FlDmPsMLF5XCv7DVM7DijaOCw8HH9+G/sxs2SuXbGI8zJtMLD9
lCiXTP64ueb81JX6kDxTXwqcm2/d6SlFQvNF68mMRfojY91rLhMmCWbDelmK2fgySatxEhjHuIoh
AXkFXbWW3QdkA6RSM25qRvwmX0OdCVue9kIihHooBDA8OinlOu7bd/Vc0U5+QNKdWdIm8UgwNKjQ
hl/bhpRsAHqOAwKnYfm9j0cRuOtdiMVIdihOreF+Bc6sTrAat20y4egsdOegwsK1q46UTPY4s119
xBhKfU9xMkOSw1Vl2HEPP4oPYvLTA25N2K1M556rTU24aXOL9no+rKC0WDXxCv3yi36vMYGJ66jT
OoULxb7xDow0Aa9N9TrDFC/taJyX70REZyodStMdcwsqYrR3F6tI+t3bvkinfmVdA5xPBiGsvyO9
LhxKxVkVui2WvA+OmWhS1muFFPB8nekXgPG905/9j3P43R+/LqzOZf0x6Fp24YhceomCvLOf2n7e
peF+PIoP9Yh0JcPzrMicB9zPB0Y1EQLuXcPLerlvkIBZkXpO2AfKZrp5yKqeTLM63bj6theyplT9
HgjsG13h1/3xUV8NCBoTdgYWIZ0unY3kKXB2huvq5CgAoT2cM5lbLOOwzGJGbyLa2Svml9+UHUSt
yAjlSjeexCIjYdnuFl0dXQMp7hBxnBU8cQe6uRIZJHp81KwlorP0NC0tNJLmRLVYhRlvpYkd6CmK
c6TL6BFHJy92oceJbVVGVcT6Hx699006N4xKMEQssVevTixgFIuSo5qIceWSifmHfzoL8pKbNs6q
AflmI7xNjd9Q4QLFt8VcFwXtinTFYhBJv/wqYX3xjfTSpNPhdaKrwsWwYECMhc/PxqoiWuXKcTn6
ospEAsOWX3l9fcBCeNj4YX1LQMv/pGi8M0cYWdTEBrlDSirjFPuKnYH0bdTGVlELfJhh4C8Yq/AO
S60qL/8xyxJTY3/CxZGqhZAXCSHn3SobpsYvPifTrCAHnjWad6fJY6WHgGdSZa4g+SZOxIZLG+1B
4TqZWINfW/CjBLRtl7BWHQfIQY/nTCDi9vgRIE8RtvlhosX3xPOXuh1KpD1HV22TzuMMHzjvTvoK
M7AwWmXB5rbTUoGEnqYAyMaY1sGOYxH0MlXTFJ7nsEbXj2tjfdLDdLQZy4UzEh7z9ju7+2ZtOcRF
kID7K/dURMhmMw9MRDvQOmKyXTbdwo8TyXrDRUDYGOAwj8pYefY8irdsyvqw4e5GlF74LEvluZzj
bISNLbOHF4LspxgH1RLunJNuJYr0r44UzN7+fvVgxIRkWoknelAhMz51g8ZIT++0rRaZxjUKJ/86
AkoQVwEnYEHx4ao8ryDGufUtiEbIyDgt3tCfdLRtUsiK83sEdJ3cMQgGXiRyZo1BgJH03TJj0mTk
ZcveCc+AQXu61n8VnkRWL/psvaS+4X4XhChXvTjJ/TseoiOwDfilk+jmo7dhnRZrDRUGVgWuWr+7
V91iCaK5iZpDrprOsf9f0btEDr4GSLSEifryrY7a7PIHB+MurpRKKgPC8wz9oTPtL32T0iekl2w6
JLWkYB9e5XcbJLo/eUpE8nweA++Atw6h8StK+7sQlERTRzTD0B8ENyP0VIayIqDdkXpBcXC4Ucw2
0tIYUv9FqwZB3VDf8SCW946Ike3n4d2HBG9OdZrc/0HER6aH14pdp19U44kzqeOaBCnycXzj//vV
BFSRk8vGHCSaLIJEvXkGQ4GDTTagW4yAThE+A5X6pby7Gg377HI7jjOIUADGuCChPj6FNjIWVPu4
J4vOHEkCorPTCLkY9Bc92EjdM0dw4RZjy3RgIiubo+j7GxXxeCpZHRvZn8oWRUuc18+Sgi7wQP55
g7/5giVOHjcxeb2VcO2fueulX3JwLp0RjIIGh3WU92lxamom7e565Yz+fnrLwd8P2gCBDmbrQ852
iVBS2IyFEDQapp4DS6UGnfDSAVhyZo+9QVn+VvmPeA1vKlP6dH7z+zNIGrWpJ8x0Qdc1aHylrvGi
isPaB9etDHYvTeWwtQXzRXeaP2OrNEcYMx6BmX6OzL8BtzKCVTYDHcGq4/8QaBsh/CV5D2HwUd41
wdh0s+bow0Kdwkmo4Pdxo3RJG8ZL0h5oY/uyw0r/IgDaH+dhAWdS1irSYwIOmMxvIrt31pLBeysW
ZW6Ikrz4gZ5/BvgtOkblSzXYVRafcXcu5TVACoMc0zrA2/4t1Uz9NdtEHZk/AWnHzj4H52Vvad7b
wbDWNHWd6eWLVGppsfWZURSmjGAqzhR/263NXwuuZ9DfKU5v09xBE7N6EnV/LS+6sEhM3kJKoB3T
0I3LIwOgVHubRo44YKyEwgJiPrbuBoKFkGlIsV5z/LcCkBq0SJ8oGgGsAWAHETUIlEtSm4KKJ7XQ
oBt5n/C0Q6Jm44Ikdm3eNHI6hDn8h8HFZhH1JVEt5xpolXofkysOqn7ZGLPiXeUW87wRIvq0nhwI
4zvuXJHcN5gyTowvuG/iBhF9QFK67HUT8ID4Vm8kXGRIUn9gFGA2Mj2aDHb1RDsKIb+3NfQp64IS
4a54IMdXJMZzHdtUvOjLU2Yxlkl/JVY8dFsMzP5GONrtSJLWQ3lwsUmGWimD2Qtv0XV0hWRteIGe
JHCfkKGBieW05P0SimXeidAnnQ5AllUthh+46FbyQ7rbMx16p4Dl7mWAL8Z4dbshepZfdQR5Uesl
fsUL/pwr9idfcCvi9bvGiPYlHJqlvpoIKlXHBAf+Vh56zEh9C4CYM5R9Lf5B8p3f0oLwD5dG93gZ
0QQ0OpcMb2YIgYclgnhSNc3iHQD5inNkDyFNJ0XQCSNuwziTH43qRssYNFRXnzwaWPBzB5a5fu/j
TpmMG8gbbd7SyUyP9dYYqAGFGXHbkbaO2icKQLZPyYTAQ9trypSJrJItGlJR/js9Y1Yvjawe+0x9
1Cyy4NxRShdmVC3uaaivuYToE7+herHKvXwXI2Qu86nlRCj34yDSz+8U2eBAoFNR0rzAeWOrDi4g
B8Wqu7VlBgXH0WiaI7oUvt+4zGG1l0SmySBAHkmJJiOaUwjHPCDNu5YwR7vUW9SqzVLzJSctHAua
OGZ8G7IBnXj1Vmz+vgMq1hzNKaFg81drSR4C/DdviP8EHznDJtMQZTRifbRUA6a3+pR5Ojc1xkfG
ZJ7WCKLvTNFbVfDXr8DQf9mUcOwiK+C2eL/3VlwT6kus46mHyiSzYOgKKoX3JfTaOvFfVEQg2d0C
SKAfCan35nOZa3Cy16kS1LkCyVfGybJw7PG7VNAbc7Nz3vVkCpQ+3HCRJ42sdAK7a14QXgmAXQSp
PTZuPwZZDcNcD+qAh7vzO3qd//Q2NcnDV/Ip/zfGEwXXGiFk57jIC/2T/u8iXPLr+oNaVp/bW1DN
Hq4+xt/wIx8/dl1s1EexZvaYjtjX+wOotKsVUQKTB1ZHBD1G13jwnjKIoSHySRj1BVoDF+x6Opn3
kk6cAbA9Ga9ZU4d1Y/obAbPWIi4+lZBz4E+mDQxKzVoxatjrsS2BhhdFT4OCZRWTvir9/44+bBhd
HQIFHSxT0DZFAG/Hk9l5a2QYtHHn37livgAlHwPj/Cgy/t5+4NvYtseJ5I4mtfVjYjzVrpohradu
+I/G8rcjFy6lUDKGzugxzO1hZqKN3VS8U8vMpzsms0a63TXpH0YPDEM6Jw90iF+ayNh/jfDNYrGy
MJuxtONmQJGNZzPhL49VUnyNgtxzrekiSdx8VxUVKy9W0t8+dbGvW46O/mkBUq15dPnxsp+PkcwZ
ehPOLb7SDFUTOaZfSvkGinHQgl15Embg4vtInqbkgbM+d54xfynEEEwBZ8Hw0U74AjnQ3KcJEI01
tSf1Lt2C0nVwLTo7uPmzDtqTpQnFFu28aG6gSVsoN6PZ3QP3mS5pOkTbZ52nOPkwNlxHKvWtKxPW
1SHb3skx5ml1rbfaLne3zPDg4lzo1TP7lyG2k6b252kwyh5WSpDopZQCHf7S8uY2aYfgo1Q2Wg32
bM9N6namjxFPddHjSF+J2vVQtNddJKsJtGNDmLAjODnxhuxmGqymYfzYPFWlOCCJfJsB+I52FtvS
TPFNJBWR9L4ECqtjRXpO2bGXGwdCKaRmZwCpD8kGLDARFqlD8La9pS/Xc8UrEg8Qja/CfLlnOWDp
n3aXuDyVVV/g5HotwiN1DnShhW5Hx+xfRt0k8eeYrX8PjHtJUyCPRSpgF3rd5Kvy3Am+J9zDqOea
ojXjUM6dXsF7fNI1MfrTqzve9pKFDDBfE/6r917A85yzvaGFJhHh90aMlGX/Ewafx0vMRA4pP96u
PLvK2AVYYJEJh/FAt0+qzIpdTMR4yxie6xU0S+fM/Ta9KIObVbkNEhNtkm3+iIpLbMZzQmcc3yGn
o9HJm7VxQgMBMXPZXvfiE6EV45gdrU7IOqkSoubP6gygpJAQmlRHw5O19958sa+wibeBqrnvEQbX
T8notRPLUw3eTwNde+K65BUDdD+Fo5bzz5FzVIaW/p6Njl9KTYd5iO1AXjiANcLrwMpU8m3aINsI
o7FmedlnzRZ2RK40QZcCbXhck/EDI2Bz/cutewBnrpXO2xEdpx1dhKiYtI6td9df2aBYv+XG/6Y0
s/0IzPKBfr9IEZA3AlrtXbhTpnHPuWaRfk8vlj6Hz2iYGE/M7hDeWyUL/j5Z//Oq3G44+za/bVSz
6e+PtBC+3T7Fb/hyPtVrKt/4B/WasgW8+Ku/1gagZz95zyaOj+HWmjr33lMsfbjfL2RTkKSjWMhE
YbLvn25qG4lYn3KKPNnDGPWQBH6TamAPeXXvhlwIhpEyGYTjpv+HzkKrW9sG/b8pJhR/2EF7AX/W
DdBcuhkivozCQufPVB7F8HHyu+oL/4kYfx0z34TOBiOgXp+WLEM4sSgyKeL7L++1qkerWWL57NWU
zFBLno3KL7RvDO1G04caXE244oFJhEBoCTux+V2reneFS6Qtb5wCj98YXTzZj1CTW4kw8CepNvdt
cuYy1ctXgawoQwQtzlFNJHIlGzJ70c+T4rSRnNFvrbsLHHaNcGTo7CnRyXOGJ+wnwR9lINXHubmN
BkUUTonHjzDR5OkLsYxPFb5126Ue/fNLtYqCSOqsQ6NFPvOs/ZaCrb3fFrLTja9srryvpClW2tqt
j6LjCWXVY5X/kkY1FePk5Y2xYpVXEZsOoBl73igHPtQt2sB8s3FKZO41CyS4GHYGNfuHOq5PPTBg
wgWKnrajRLY2bHpeTattoaLytx8jMLg37sGlR3cGBXs9TTX7WRwDAXluIHi7L7AuWKrmRoh9TjIR
z419ZRKwbtnmq4vSSXG46XJKZZHMmHiMYklEx0vBSBeC/pdc4VPvkU8idbkeM6ez5UQvGB3d5sL0
C+74S7CUqHVZGF0Z4kJJFFpNhrs5tC624/fiaOj54U3HIFYeGZGwlBAcvp9mXxSUApAm0h8Waa7o
+je5UK8spwOEoaQ3h4gQzrsOSrmHb3pLRnr4MGgIZ3MIoJP/e/6QMFp7DJfgo7Gw5blrxDeSD9io
Z8MYL0/sjNBLLUooojsMP8kshsaOd1Hb6Ml7Z5rdF6VlNBRw9v2i4Syy8Sc5048Kh9zpZBq9irQb
CeVvrbYp6r9rfEDOuVD9yW+Iku5HJ46oN3/r/pxJXc6Lw0vMehZH2EOPl0HVcKEgs9Scy29BVm56
xGUc8v+SOnnFAUQ04Bq5zrBzq58eDQVp0zMzH82ab+xADG+QM0ezQ09xAl3/bQUnLDcNel4bn1WT
zlUDvzzNEEW6arF8TgZutdXygm1ni5Wa+B+lDt5Ktk6XpijCZ4IeDWPyUAWQ9yKSM7N7k4q9ymt+
CpcJXta9DM/FLyJmrbMnWsW5plAIaDT9naFqb2UYG+t9EfUJV9kC97AkBRQK1NrNqm55cfNY0NG3
WAbX5UmRqey6M7snsE9iDmi5yfTZbcd3jQ360OON7Vrxj9VVov5+zDpjsVnKRyzr2tLPA/4YAR2D
Nxa5GXHtDKFAR0V1N7oBlR1VnkGz2mieRI5gcgnJpEQ2028FdxCrvz/FyHsyk66RLxJlS1KdyR7D
LfHe0Yu824Zj6ycdvmysXWH7OUINgGiAV/QLuSqimJBvyrTo+xVa4LAF++Y+6GPKqd1GS7pKP9hj
vkaL6OPQfpwiuuYxrvtpq1jPvgtcT4goAI8d01yRVaH5eYXBMMyzQ5DERRZ/H31fSF2qYWu/r7PW
6+WVhtc+pocQcq+EfoAg8UDoNmMg4d2OWtJsGuTFlRVhIoa8oHymAQJ0CwUX9k6FFMqmBy8tTH2z
2mIqxOXWbZg9LIufUCHErWh0GmBZNK1xaTjP37bVkoqrQNdWmx1XSRco1aTAySAvjzXdYnd9627b
UIYu6pGSQTY7Wyh5oYGBtpHeru3NwHt4VVwvBc+/ASGPB/rr9fACD4KpspvqnQa8SjnbC7DUlRT4
wPJ5VlL8jhetnHnvl9ZaCTVsOizcrWH5Ymc4eSU34wz/sH4XVuHE75FfQBEzKkJbKR8ee2yoybMA
Pp8+stnr4A3oY0sCu6D7CKAU1gyBAdZ0o5rjDTfLTiQOWiSewL18xcqB/YslH2fEKmW96tld8PfA
BM8p0ip4ITbkpzfK2OOEUmiSpQcbaTbZag1WduokZh6oAEroNq9VDTFI07imAhi7rOdj1JUrYAks
6DUV69lfaJluXuBCE4sk/Y+c6untdoxOadZPDfTd9uOl5qmiCr9+jAVhndo2udziqu780eqvs/37
hgfzg0sgV0uW5nDgN/9G2aHGLGauWSHlVhgzLpfp7OLmYB9u6TO5WUB3OEUnQ8UulUPj8DJCGZFN
Bwk87sqJDEwYnfVKvkin6fiYDhKQ5SiYJBgODSH/n2fSX373eR/SLlY48o7zJE8IZnWQqBMHz2T7
s2FiqknM72ahNWhgEfaTk+N/cL1Vp02U1tXFgceGx2ogJl2f00s9HTbpHMs89pjJt/xP4zHCXBga
x+yppkOnyP5/mi2seDskz4gmIqEbxLCo5vxIlgb9dVxPjqzF+sTfLyc8ySrO0bvEgmjZGpP3BDqF
TPmglZUUNT4O+LblyyCVsK58QJoR8WIDDGLdG6U9acTLBjAI6i1I8pBRaMx4ivmjUB3Ucmxj1emz
0Y3xBIaYAC3Az8TG4f/S3jMDAaX0V7jthdbNF4IsDAUUiwwopbSCYDxOju36MLVIvPTEgUsc8Ocs
3kZT5z+E6+t308BUSvpt5hMNQCi6AHfzFF5rLUpl9gQh1a2uPsTuS+eFZfZkUZDLi7ANqAQDBYw1
39Lh/RD8k/QVDHjaNVc/LxOVl18qefQOKjYHk6/bZK8yLWQxl+epQIuFQvbvcidHnS7IhmaLqI1Z
fzRp2NfQTLBBAsP7gCBgsFIhxbRBGaJkwdDVDVU/bE0uHkAyh8XTTE6QVoS5sgehsRr9mM9njinz
UJbr2p8OhKtPi2iD5XiUbv9ovHwo60SHeuOoTXI696PV9laSxL20wfzjXMKz1elTTi2Cuwxi3KCA
HjxWVNgKC6Jz/WGSgAFK3GhpDauNQeUPSuK5sDGBESPVR5/pgplGKSlEBgRfv+gLZKcVdUbEk9RF
Vl/UC6Nref0ol7SjnUzf7MxwwLCVH8PchaqMyjq6NF14a5iJNoA19NmcxqXRwIXVe8h/r6fhU2iw
wuX3ktOZ4HIFxOVwldRMqOeHMmFuaz3DhK4Eyg7nlvVcWB8zCf76R7j2hwJ/4SLqsI2ccWjQUngi
aRokRvwTi7RnhZpbnDI5RdQpiEeOv+AUxP9+9MIP5P4cyxnapou96rDz4wCnHl2lqXvUxLn8N7Lt
4hkhBNt9ejnnOl55odWBz81DiFYUdBFvGEkq8eIE3BIsg746EvFSZUKuJVXpFfLvlxKzJGgXjn0N
sP3tsklWB3TRp29lEwZVJD4paYU/YkRQMjPGSkRzfSpx9dGL8zeXNJM1ACWjl8erzmolN1R60Iqs
J3dB5cqsy+61dYdfiF2Y/3WXmuoGrHFXg36VrWxVLFmePjMzzHKI5GRPNw2wX3cy42tE8XL10nU/
iqh2hTkgQ8FBQj0VjZZW716eHzwBsI/2NN9o+R+8BBlVEUymaqcL99+P4B03yIlEyq6AcSQPSsb7
TGTdJYHzk4MU+737+m+mDpD1nIYNjx2rX/ltLuADkD5EZEhc6gF78wVbmU9KyVPNaoVyJMlGlTsC
LfgW9/O49BFGGlPADei9MsmWFkt2b2N+A1Vakr4vBGHACBDj22HsAtwKegc7MuOdrPxDnrPmHe9a
swRfmjFGfqaNaYgBy4IEZpqCTqdu+0SUrNzGF/n43cNa7E0s65gt9Jn1j05nXZ3xCJzsfE0uwtPd
ji9TklPANcO0RYsqLzc45ZTA7+NlsNpdbjDf/WEQzq2xcyRnhEWTKIWeRGThDON9iFPVTP1JALzg
Q/CE2i1hQK4uRuoCVNkXOAskkhipv/kz2ZKehoNM9mO40KzfyONA1voFUrW1Yu/BsDmtE0mPpmX/
UpYUNdJX/V8ZajIRHVu87ydy+qEHCNGtEtBPZM9xzFtDozSoHUn97cM90UKzpDw5UZ3MysgfsPPO
zYhw5SraIQI4A/0Z0yZk8OtOk/dSQkwPcsGBhTAIQ/cKrpFXRKYOWmM6ekUlXbAdw6aP22H6v1yD
7FbaYq1FWhaWnGX8NSS1AUjcSXcHEuUEfJh5yCEnoAQhDTt9vTD6s5E3/zXShOHws8l/ntjEv3B4
W+myXJNkAp8hKZWpoyEy54Of6U5x1b8TuZjWnO0LYyF1YOH6UFfVUMM+uGo2YABDyHr+q962ZAjV
hd4RN8PqY9roB5Nh1cf/f/fPOXOPQqzOaL66Nd2tyMdxw6m6HQvhBxuRCvBQgXfuAiRm6Gu2zKOd
1hvzV82eGS3G5ks/VRpqNhba7R2M+Y8+lVrLXVIgwSgo0C7vNXZA5qp5YCaqbUK+V7MUmDP5CyCU
JIJVya3zxhMnXuLlLWxy9Xl6Ie+6t9jjd3BrEM16FYVfdxwQzdF23jtay+BXjxMzFEAWEAydCCIA
G+ysIW8RBhIx1cLwJeaZScpd8I+NBPp7Uu8cwR0kdwQUahia4+EWYqP47W/f02GAEFNXlnUVmI6e
26SI5DXIfULZ85+OXS0KT+6qzHoYD8BT9E6ipdKOiGzFygNlusnJCTx+y4Cn8SE3DteoyiQtGUK9
z4PevnXgixnDQqoffK64c2jOs3GvO+HiA2JqCcYRzylIKnZZ+xvIshTct/6rCG7yszfRF+17DpEo
V99BhGOigZrYqm8zX+GqgfF1zfrU3F3UUxDHtjBVrWJm+zZeGSVFCToW/sSLUWbYqnwKlACnLkqX
KwwRcGowL7LNJjpD9AdiskR0UhP6qhqjFmXFRgaRAqQd97CnCMSrrwisRAwOS3bMhbQhQ+Uv//0v
e3WxBClgvMSSJk0bXKlMZ+gFHKmbx57PktEKLYd24se6nqymw3t8ybayfNkNMkBeQYucfFdIaJl2
WHAf9/p53eDYp4CY6sZe0KhZl+cvzzCLkZ+z9OicNZlctj0KULUPXBKFew5/tXeUy7gK6npQqWWp
M7MZ8OIetZ/Y2wcl4Ioo7Zbq1yQdm7kyqe6dQDWGlw2LAAPBU33UrTb+wzEoW5JfpLzoyGyhb0WO
0uFV5+AuCp8+UCsfJ/ksDL4LX+Mp68DA7f0cQRyQbD6/IFkvGfyiHCcmxdK1LzpHdhoId9RchBkk
5nawiSW4R1FneG/3S1P3pdK4I7SvnKrnjXtonp0RMBEM7qkXoOVqhHM9eQN5QXpdNspZd6/pUUpX
vNWvGD7Q/wxj4Fi1LnbBAp9H/J7DS3V9KTiT1lY2taCbyHgrrZdlC0LYgesTSTSsy07weYQIsAZu
Qa9Iw3Hdkp0PEVNtqLr2rk+ewGWlFbBgfNDZKHgd6QAZsImq9ZMcRSne0igwy3MrUkXGTC1y81kv
OKNuMg0eMo/HfLblTspxJJzfKW7HCggqEzjqaO7dNA3S0U52nXfTbgWEZAb/QiGA/kAMdp5Pueg1
p+08Ew4RVFrsFL8wQc5Rp2qnbRecVsnZaPOBpWkpnam5wEpbDQRe6j6Ev7sONARa46kwmtHsMjkI
0uDaDac6HXACIGfkgHAuOaNremmwPXc44o07RhePzZEKLKK2OOl9Pr7uRIaLkTKrNQ8OrPSAgSlD
Fsm4FBtNh5kPaOOSNRGMIlJtg3/UkvFdu8/wOyDPhJ+wBpKwKMkeKGV/GbXWc5Q9Au+ZOT3Ghvko
PLJmTKKgvsxLQJebm1hgPPMLcyYYEakHnqh34q7smF/EJgtWYXlvoSgPKl0MCVuGNRso0fmeJeK3
Q9V4o35Ekk4GUyFoTLSKYyGH1eOmGlcHhr7LuMTWlC3iPkfSrTIxZs9aSBz6sB8JMKL01+cIaby0
u9irTF1nDh4y92dxuFv4rfNMVySQ29hs9+9jlbXGq/5qFTh8cPJNBrIZU5sFus0oPsiniRtg+PkO
+rO3d5fvCSfn6IeOdN4VhN1VlnPza1zO2dem2Vy687r7/POljjhnhw5mpawJYAPmeavGdD/EwbzP
AyREWbWvaY788dllza7O4YAFVLqFXOTssxQ9VOL2yZlzcEXtMoJIgA9uI+/fqTEzKZnuMZOcZVNP
k0T5/gBdIjW/cu6EMG/6cH7yAoz/LcvFJIZ0e8Q2ByxQNiuE8Qqf0L7sCaz7jk8AoYM4sLNNwaGk
NOeEcH6/ic7TESpLrjPTqAkShEwYcV0LZTxtjylAI2uJVtIPEuI/6Gx6VB/gyIRbn5wl2qW4LcMZ
VqfuRpkB0/AkNopcmv1BvnmUFOriqx1/LJublDgiK0G5jI6iqzgGQUETZLQoXJBT7DiDjzzoy3b0
ELapsht6VUDpZBtkCIenud4ZcpJWygTXcyFETa4beSP5RmwSGi8C1WzrEcqZiUt7afEtQpQaIp2z
HbGoaEjNhkiHGyTHFtZKlXyu7/pMhnWWgHJjhWbUI8FAaP3916cHrM4ju/VxmXnYl4k/b6gk/rv9
JTXLPwVu9hiYw4zDkK11tmis9XITWYrni8Mmk0dUGkSYe3YgOeg3nPD9/hMA5d+YIJRFZNUUDOxP
1lxVlnH+L76/Mn0YGFTEbn0aqxTsFM1CK5yGIgQcwFus0I3SZHyVK7f8zHXsHWkLe2GtBF2yipnU
Gt00zfW/IdDw0Rs+G4TjbZJaJrCRy1vPl9HkK3ctuMvFAbYESQ9U9vZi5298hfKUKGuOelwiH4lf
j6pqzCP+5PFdp5AMWZKcqHlD215eNYK+YyH3sFhUy6YB/KTPN2xhmAld4H2T1tYmlYWTHS7xPgvk
f5hlvl4HiCJAW7NV9suYAZEqDJYHbsru8tYdrlawmg9suMVpxlOdLmhdjqs+CNu+bgRHo7GdlaIh
hCaOCBhrLVXzwwG7buO3z0rCsv2aaGztsDHRb+VcWPmttCFf4Jxopx8yjCGN69AfP2Y906eOkRpb
1/CpawMOQWg4sy44tWDGBf1qd4vdJwwClkuBb1WHAGXx7bSknRMy4XKK49OsL4if+Tq3zLsZd00D
jY91G2BwMGxpQCDg9HWkK64OOYzjUdtPmtHUELkdxQf6deMcvPsdOaaaSaGwQKH2lH23DY4baQAE
pryqNduyQnBjWw1aFZjhpZe9m0KGsdWbEaZyY7Wtjtl47PHOQoZc6VMIqXslUeGmrzPALZUYUWCN
MvP7+d2+nlkSXkgbxNZKwygtleqh58OExhme8ZcE4iUC8R3ikT7LRIV6ffIP3xiEbtGPD0Ek7g+b
fUCMozwFBHCzh85S27Y9Nmj8tOe3xrXOyjFu/Mmntim72iaURh8KJI0aXpYVXYZ4rrN1ARNl8ArJ
divLXJm5g9iSP3V93PXr52Fav7BZopBE7ildQhZ7KLykuD9H9mquV3afP+CxAHxb7spUxdZnRmFE
SyOL8IZ10TzPx6AdKfSwBqtPD4X9PHbj525JsLuibQZJW0yYtVt0CkFwhd9KFd2urfzKYRPdw+QJ
Fc8XfGXlG6zg2wHftUcj79/6eXMUPkUmZc8Kz1YNKJrtbB1ArktSnkzcVVNLFPU1/kkl1RtR3f62
g5u2I5bznJG+KeTce8PDmsZICkPmVUMC5d80oi3/jR21Pw1WYA+tUnQ6CFCC/kT926pcwf6LBmoL
qQMlh4uymXtWneAJG/porTiLD3Cp/XvZ4byQbdBUEKNXDF70+yztwo/p3YM1axNL0g06d21V5W0y
eBRLjfq5ftakUa3KUhMltMcfQAeQrb0MNXNxNmT7lgYbuexU07M56r/7/RVOHFfTjCKZTXcW09X2
Oxl1r7MEIV7F4HtwwXl1DY978xCgZs5wR/L3R/zDnFDgvAfyMT3Iwp/HW+6uPtzxG+HX6E1YsGDk
loNHXlJkbyVtVuZGZM/QtkE3BzLcl5rRrisIE5rvaMWVq63uC0ea8NnVcnq9WW81UrwM0e/ZGtnK
jzQ6eSdMJ95s8tXkm2ui8poTw6duCfCLtYC+USDDphOb6UmBq0PDfi5YrtEMpO9VYQ7Cf0/nlw+i
zfopqzwRtk3rNnbxaetFNsgIanV+it3dBCoU4mAe6p0EhHrpm0OBNL3eYMvNQhDfluQhXsyNxXzI
rIiTWU3uIVNnSzzIyXn/TRYm1BVDoGaPI/lBj9+0QzMSfr/Op2AetWevpwch7EdRrUljG7t79x/8
C+IvGGT53xHu2P6yFQySD4S8i5zftz5RLKsg418fnoArCjPwTU94CrVDCbakbz/CAWIHDRW5Rmve
KSjxk7GfXBbthjOd8tVkxPrprdtmQTuQtkE5Rwx6yMdHgSbSecVW1WYZcXe+zJh73YoN4L1YTzry
U7MMc7a5cA+St3PFYF/w/qU1xnpHmRL3tKKv830q7lxpD4VLT6WWF8HS6krkrjMSFFAg3wZ3M2Zi
GcFdRGCS9zHHBoCi4JBusUBN0bFXbr35Lb4LX7TDpmtv0cWVO/BdWVkQNh28xn2EA4jSmWcZH+j4
c0Jy1SNrP/+xVY1Dwfo2AyXHkeA93i47J8vIEtVYnyU6Q3C6JR8PIv4kiBk/6Ml1VcuvPOO0ApHV
OjCc9jM0CtJXAAJu6tfGAEETBFzvQAJtfPKNElaFNESi2K34qgoI0cbXeZMg4NaVbsA8ul4roipW
7kM+8okViCCzxNIQ01FpUjPAj9y/T9fEy3jLB1/SbIo3T3gOyxjkDkc8QmsUwgNtYidii3dI4CwS
Yd2GIJbiCKr3rBJ/P9DnTQku4jyn3ss5aON1CgHcgooyVGcxyMKKbR7N9c1Dkn40ia2Y55ylzR7+
OFZDEBobKHhiCcvHuIY5jRUoDPk9FapRwW6u1ANk7htAE7Ke3yJyeiVYrV3kWkpeReBba0Fg0CMH
t4YrX4iQLyzDTs9I4JiF4ANL2/Ms3EmogTf3m31AsUWwpwRRAsvuHyG2H7i0SOMSZxlFC8R/E+0d
QxS6LN4u6tWZ3rdQoTTzSgxbwpxgrEBqK7ykuZ++aALXhEL4nRD35t6gmrpxOmK22NpEARrT539r
1d1FFyq2lj8U+nGyS30TAFcwsM/K8RpkqcqiVvTZjNxZR4uA9W/4N/dyo8GOjZ/IjW17QLSbS/uI
J57EXKWPqHzIZ+6T2gz/ETSr29ocO0QyTpWlvAEb9HGm5DJ2dUdwlWw+5dPiIF/Mbmj/XjVaMcZf
2Kg4EzYoQbKsSqoLZ7GeD2a2Q/nW1jJzB+Kw3MirI1OVxNjx4hBfhde5rHUpwexta0xQtEj4SmQ/
YQonOFgjmSxW12++smIWgM29kQaUniJTeqj3O2FH2y6QThPN9qdcnTHY5JTGEhGMZlPEQ1+aaRsC
uVJ7ugu+pnvrrsLLlb3IMLi0NvyAPbvBpEqdX1QnXPUz1+RmDOozsMG4WMo/mQtG3CaQ+/YRKkO6
MW+LUr8Chy6aAOLY1kgpkLAyKt2ibthfIpzJfEctUtWk101kANN6+yAxi0dZf5b5z31+aCaicUDW
gccINbB0zS/2elb3obqgIgGWRUygEYrjQZuL48n3S21GYnTpkzIvHKe/0X555EEknJGnDKtNVUgh
re6NOJ9uUZ0wdnCVNUvHKi0AykGWZjXjbVxug28nCj5nvu1jL9cqz01oPC5PGD11By0QSUFwnyC/
QcTO88sbeIJorZEziw49w/dShrA2FgtlC7czQEarDk9ydJPHCKYZ+A8cJVEeYUOyv1hTVw4yaqvE
oNAxHGn6WrgbD+GEwItc7kl4kajDepgTo8S95nTP3WSB63prvmOWCKV0qNrp+moI49IilafQna94
73GdrdO0BlhO6hnYXZ792CwSeovRtWkL5KQ0UHUlK+UpnRFWqNRHWaUcafZ4ujCGYUtbVD/X8ycg
tlM/DobSYxtYAd/tNhFg8SkaWVjSU9SZ5Av51CZfGRijRMAIpjlV8dE9X9tv5TyJ/pfdWxkzSfdU
rhMzGqCob1UUPBy5MsCt81CiBjfQ0Za8QqbVo+S0rW3dNzObkT2e7xCZlLUfQ3D8EkJldzo56QKe
6HsTS5+bIlFiP1gey/L3pEx6vTm+D1DmytGhTnjmU9KJePFPFN+NOXlkT8RIOUtOWj4PxcmrXtzT
ksItZ2VyF3a20cmq/ZsJ+BbkcPSMb6HQAnzO6ADsvnridUhgmrAFqmjEEwvhLVcfGXWOFUxDYdOm
tNynr9WWHbz6HYkZc1r/1oXXXNZiu6AtFIIcIyhH3SJ0Igrgqy9aXUCctooc2fiw3WIbyqrDLPx8
MVQdWoboZIHznyxCRoUtPFN5pWxrQVplcm2XjNB07eoWqLnFvM04TzM9H70/jPS+GVwH6DMH7Mbr
Dhicp3a0OdzDKgb0UyCVkNnzsHowxYxzjDQkgESN3MIn5fA0vtNsRXpTf7SiJblKvcF4tLIso8pG
yT5YYJWya7v0WR9Emp78EOS3QgDQZgj+p8MyFoMIPrHNw3x1F53dtrK43XZc35kaTzSTsNLsBMxM
91abVQuWR39WOisALn9h1txjWmT71GQULR7sXP0inaLCMC1jmJAtnvdgzqwszfqvG/ksrKul7u6q
JPWIzQz3N3JC5rEROIWnzxwr4dmo1PijdeJHnusAxXG/fZ7dzMEzXeCGLFQMRtXIz1/xuLT/q19C
+HazAukeiB1uv76nDSBslRYU6KUI75zwXPp0pQO16O6zhaXWVRgD1H0FMNISivEmZTlrrOv71cx9
14A7bdMfTv+zMQQf0hBoDy1CliU3DTCzbrpEWKPw4buGcR7BxqqSs3N97DXjtfCLf5DYyvzM3gk/
lzwiL+h3uRxdWVN1JyinPpOTuWKPZ9u55FsMOfbBZDEk0ck+EmRnEEUdD0iyFV2EcCwMzBjfo5XP
MUP0cHM2oAtT/qM6YammoJVQb59vkGWjSEBK7OhvsJJr/c4OOA8dYMMIqAceNz4yCtSbCqk2Wnyi
r9gem+l8Rgx0lPl3hz2e3+GMfghIFDbmh/2YLl6b6hrNWncjZVtgg9rXM5ziEXlE6oiLKPd/d5ou
1CfpP/kvsjgLIfgRZhD1gQ27HEcKlhkLMEi8zq0TlE2zStnvsEPBpfJuLg9BiNp4rM4x9QGkAhin
3IUD9T4YrUCl0Z2yoelmlyZIJopYnAg4zKxBQzJNwX7xhxYuwQZv4avdhcHVimWqrjoL6LUCJDie
HQL25pqri6FrxKcUcB5xZmTa7w/qUUkgbbR+edRrtcVh4SR3LEptWG6tyaR2AZbwSs7ufd4p9pD2
XmayTWm+ldfBJGwzckNwrWwIGXwOt2p6PI6FoNj1yAvDW7w8nu1RqCp+QxHCF6O7n+gDNfD/0w4R
GUMHCLOmSplnKORAQxWJjm2ueSrFuYoTxYQP/2LuRFTf/FOkbqjG7Yfv4FGP/rS3WfUevfVmGNDg
3OVBNbEH1Jm6c/PpBHuK+XvVCw2AHzTMAtKOEouJOxJ6rqqbJg1QxfDV8lavkjuEcDVbIa/6QPwx
qpr5/5AJI9DyMeIM6ZhZh+lZr+6WP1gUPZnJeRgvTrxtCvykMOy0HE2DO5uHuCoapo4K6UJYdPIq
6u9rkctLnaN2B5D0g+o9rD4w3cyE6BCMJa35lSgSs8kpzzZ6fspfxc3HY34mBwz9BVJWIyBLwI+2
RPPXeaEVvstOpdL0zwnoVw0mSjH6AyS4W8kM4NcWQnE2YfMNgW+Td913qA7iCvV5+nzlbp/5igBA
wQ0Bwq3uYTImdcc8M9ZBkJSaP9y4S0N7mqQ17x9JnsqWl5gHy12APoqvykV4KZEovDcJ4l8Gd43R
joE57KT1KO8RBj0Dw6ob2ZMyjb/YeCymr6gGb7jTAl+kXmpXzXytUaybbhLGt42D7+FfBSa4mRvj
kPCGW19vK50lZzv02ccSZSEqIMxGjGVVBQxowJYFQF+0HoEFX2RObJYNz4D6sOh1asHvZJydw+R5
pmMjGlZT2xd3VWyRDwA6RfQB/qBtfEIaY4ibXzu0wLHKxK+Az1CfnwbCWBZSlwjShWysFHQOBAJf
Clxw8+PGtbrAtt/m50eAlDs3i3+ZW/sd6wQuO6SKdp8xUG7w4Hi1iQVFzZOpYDESvVXXWC7D+hAz
Ch81mwwri101qWGt6p0qa2sBd7q6fOrcEBRe1UJnwqsXlEDjRHn83AENYC99wot7OoLENiWDMfx3
c3rlmBRnUI6tvzphTT3oqDAUPGPzh/8AxeN63PJmyxtzNv7jwJi54hbkZK35WZBd7aI/3ug8P1P8
NPPxvbR39P5Q1tkD+I4l/6Tl7tWpo2gKSBQHjF6+R/bHlUU28qdJjiS6cSnP97edZsjv+87dfV/l
v1xmT5eCuas2JH7V5GxUT24oZwn9o99cO7q+qH/CVF1VKr67JADikFjDGmb+0v87AP/2GvL1PV64
oxdZVFo56JVFGcb5b5l12+a4x1dFLP/GxzDcl9jZvc55aWKK8fwmoeFx7ZKYA8J9BgAOEpQefYec
4qedZc5/i07AM88xzrvzuLsufl+mTcAwAZEKe2qKTbSt7+TUMs2sl95eKjNswLU7qZETWMTs6ixG
XL8DPoQkZ4qeMeL2wa/zL5rrC1QtmGckJ4eWUKRADHeQTMASKNDFE5Y9P2+EN1GWlM0JrleJchvv
r6xRcxJt/AXNhbB6+Ow6JyB8iHgBhvTBLq7U3BMtMwmiBi2rDEFFN7zBlahynyDK93rAJSHXIQK4
CI2gOSelj5Eq6WAd3JTU6ftmymLh7lH3ayTCCnFO7iz7+uV0XcoDSvzBnKK+arh/A01ewUhlJIk2
6a0PhuzDt6LfEB5XJNBJJtVMMH2I8Vg5b5QmIJogTKLJgSvpuzZOIbZQnEDn/IoSfOud3y9BdDDL
tqhjPpl2yFdb00vZRuZblY4Ow0pyYV78BOxbo92Ifh04cctP2xh0mYP+W4nIMIpmKUga1JWMrCdf
8G0w3b7D+AjTbhB6yg9JHrlcX70hwPuNpRRulRUHuDqgqihrcL3YyjPXzO2zZK64i0D/vkQ7gjV8
4NYMFMhh8CVRZoGiM5BFtfKHQ8i0A5ju1wjQxTT9xRaSDW+cUWFycxSJ15+NXntbL2HXAqBm2aBQ
VjVUCyXP+8p8on5501/My1hoOv+Ke16sJYZo6X5axip+ZAjaiiG9IfVMmq9iOWA3YunP0K2qbA9U
5h8s+2rNFaOFAFPhSEGkkXM8/78L6uhIjqHoW+j8rntIvv5ID7S4J1tTbKWkAwwnRlqgalhWe3jD
RE4dfHsHTD/I/YBCIP6enyhBIsTd3j3YoIraejMfGOo+LeWIsWFCrtVFUZaQRvzkGfSL8jOik2Ig
r+Rw8das/ox8j3hf2yh7xdG16nUCZU7YAKCdRwGGcDMN0+PLxrdqzeUbhsIRrvyQls2K3BLeHnWy
/cfKVlqrxTPXypw6Npyn+6z809FH3BPVtYwJ5JCk/W51OBZcn+WM4ULVvwgbTUWr5AoD3N10soNy
BUbguGtPHn5QITaqOGzk6EkzYq9ZjE8U7OlhQrhsm4ilu9J5DCUzCQQ8dBhOcB1AVmFQ2rE74lcb
2Zfhrf7qytMr9A7VdR/YKBVxztqq7eHEUWkHJlplGP7/+nvHgNAB1iLF1s2ZxowesVi51aOXP/l3
lY7ir7yX3JFOhbr5dMZx8HdHmcMCvM3E+bkhEusvms+j6bq3Ab/2KQg0dmt1rNizaO7WBP8F7PDE
Lmo0b2dNGZU1tuRe3MnE1T6TkEzcVaDfCFPGlPscx4NIhhogBV8zjW0uxaTazdt3f5CTJg6NWA2L
M2KbBVhUdH/ud/Ioht5oyYzAD+yKbHHQgB1tb66lCweuT6oPEVTlfhfOZY+nwzfqVdcMy4aqtpzP
aq3WhMqNEcirnP2kkd1qS39gn1XUbwIVkUsDfYA+xGzwecA1iQtPsbvgzVOl1jzd2FqpzHONjcWx
wEvLyOuWt1hFSRrWI5FW2ggDxY9oJmG+rxISoosIJM5EQtBbnddjwrJviHj441Pvl761K+tBIYJx
1mdeYYj93v0vekervm+SlWshxOqTUrrkuhUMjp5IlOWfDJ3OS/J5AL+N9MPWFlKMH3clSsPacDZ7
GXVcymP3znnNAI9EoLOXH8Kcg6nAHIYfWAExTOtRDICalS+bnTeX5RNjiBxHf1t4Xw97/kwCmZh2
6f1vkcebqwnwgjiQ6m9khNHDPWxYjtEnEh0StvjOtIWBgmk1X9+wFgDNy+YU6UyQAwT0l3Z8lI7V
UQfS6disIc5cO7SxeQ6qrbO8Wqdb5D8rdA6t8UPM+rk9+Fot1pHlOwEiqNdCQW3iRnxtrBTa0o47
ptvzF2gtdisstNXsM+EnNjy0oh/x8X7QPDQFkYb7tA9tmGdVWS/djhsrRU1MlKorcW152D9DCEN3
KqiJ2ntPDif4y452qSB0UGwOQhUfpVXxqLfRl7Bj1amyYFLewW/NGxOd/1AQ4kaHn4q7pr3xC1Bl
NBSDeD8yDVAhZrt1dAdZo1Xu/yNS3UcmjsY4EksTmqCRH+OROz2DZ9QxKVgzBAAlZN7CXanHZzFM
sE8ANH75EcjGwWG3co76dCXqC1ATrt9gE9dwp60Y0EALqdTJC+Xv23TKlJW7JNxzgMoOafdWstyF
wMgf0PoWY0vmql3Q7TvBBqxwrczl47q874GCH6IRtuNxv09sf1RVryai3U0JWxOOke2O6PJkGl9J
mdmjLMqWFaYjyDwC5riq6bi/gQ1Nki70pGPIt5ovZI4ZElGyPbh1L7LOOCpzhcKDsJDscHjdmxnY
TiTz8Pi0uapgv4QUqc1bn+MR0Nz+W4uYCZkiH0L9wj/EF9aMpBMqO02aEFlM93diFVAksNbiatRS
18HURl+JVzvw2RCeA1twwpMzZgKCZ7UGrHFBgFR2DvZkpifpM2hYLjHrHICBLSKFKVwI8JqUUmpS
ObRLDPwfDe9Y695zioDo3LDljVfdC2yk7GBIIIKM4bKID8PslQUtCmFJB44VDye8GiY0wvWMsDj/
w1IUXlh0mygRGhnJGbn+QGMOnCAtUkRfHQQKoGVdCczdHm6TdVTO9qDPMaBG+e72Z95h0U59JNut
4PxNkEQ/2vMRcHTCa0pzUTliQngvLuenUfhiVtHH/21TTCYpf3Ym92rHkdL23j6VG7GxgbHvmQfa
+3FDG1Evt2yhyb4ikTn8hGn3+d5tLZXxK84HyzKLFiu0ka1MpRXyNmhHVSk6BXc0Ec56g6Cs7AVk
uGUHb4y5zbMql/W0/bHF7PR6tR63wLtcic7kLrzOt8OEMnOGl1CVZwOfq7zX/tQuFSn4WZXFPD6G
SrS8aSbV62jkWkAO6JjGWHT6xn6jqbsiptmJRjaRWpvzs5x05p+f+6dteh9CVSBHpKLy8302itH0
e27/K3veOx/lzE+3njbbqiTQOeFn8Fnm9RORoEUqzwtlZ1YCldyA5JhlCbWYWmdNFSnqOcgMO49C
UWj52xuYnEwz1wFSvqDLYfN12/TS2ZswZ8uopJUktW4+5iq43dpOtepoFVhSB0TCnO9P8Ok5hUV9
/rdhq/X7l40vqSXRP/usEJTv9ugJSDAJlC0LBMo7J9QP4OWpq4t7Qu412AEPhvgCaai7NRznnyJV
TLW/zMZ0P8rPi/xh16rRvNL6uQfxgUf97xGSUn9PX/UMcnGAukUQC2SM/TL6zzUvqEdoC7mYWBZ5
OvtI+w73lQ6OaiXtImhAmUjpFAlMO0iP5+tEGDdWOnY6jzpsfkB50gX74GUr08Lf2HnBBUkOyF92
D70VpbiWyzrQl6WRBa6nKcrG/ZJx4ra80zCpC/UlFFeJYWYo6efvvkUMmZOeVsiTguvTefIJWL4Y
p/5Aja8pjKmnJcN2W1LeD/zmPbP/JWHK5rbnKJ+Wl5rGBwHL+0nuXRImyHtkdhDnTceWwNK/suWR
S9kpyyP4DRtZs/lFx9f7mayjKx1l9uELqADiT0mt9qJtEyRf9whayLyN22W52mOpPRNujVvjuBxe
9ekT43zjiz6cm7rTCml7usvmik1L5HSuVmRyktGDjr/w4+7UMT2ZarJLKeolUhqUZ47EXvc3bdhG
XRUl5Mi4QyZgBhkk7hgsrHsTlWKtQrL4v84dQa1PH4DpPyagbCmi525oO6CTnuteIdAkoEeBMp39
oYyTbAZUm4dXcdr2fZyOJ07yyKvQfz5GbBPXidDYWP55I2JEVz26hmTsJCLzT2m5a9w0WU3Il4wL
7rVrc7bPe+fDnjQ3u71/DjZaanPOlK/lT3VAIs2FTG95jVzrSjNhLA7CTqza5ahn2wWS3ZRhiZXk
/qpix7m/9ZazqaDim/vqJLMHnmygvJPk9id/PYwRosHBNjQLyRygc7LcQBTW+oipTkgnCEKS8ABO
d3F4zmWssdJhmoNh9QVZ5M2VjVlx19sx5ekr0UXmL9e30L/ebzEeJ9ZIj4UA9VlVwshfU9oADVCa
kvI2lid2XIr3lS7q9WAR5Cb9bL4MZf9NFxNsO5QHjgkMiLhLgkYVOsd8iFWcmDZ4SAq4H4Ii90iB
ks1V356DuNZTZe7Q2lrWaG6ojE1G99BQUBBapTNFxWoMjgVoIhd3M68oGySF3dl8kMk5e2on4qnn
KXKAwka88gwc6+Rk2Uilv+VBB8bjeBn2bB7aSXnCA9WCuB+uy+dA4qh9C3cT2GJkWxrCYyagu90D
cB00JgXkXA+B2NqQGEdgNuA7wOo+Q7dTShM5HW4v+fDIoe+n3r6M6TnHnSnVVTICPsESs25hu5Kt
x/A79tkTE9/cC951mbtC9XnYkifaXR03554YZpwtFhIZOCNLpGWNTxGYFjr+M1bVb//IiHljNS6F
QAXiE59CNgjjG6xwKcYRRig5o5YvefpYv+jdfwDl6In2rnwQz4OUobbQta5aT05b9osaBbI/OyGU
gCqbvmAU5WbMAdeka47WvImuEQmUyiQ81y+XdWFHDX3h0/co60G5WFtWMRw4bERD16BCGAolsfBS
yLN44Gl1jgP9dOlSDbBUZnlx2CUexhpRItEFsjUS6StRoIRhhHulrVa3bnHrztV2dOab0JqfLhEs
PVaXSj8tsPZFGMShlxU57FhbdLjBB2c9/Gu/plKsBGEgJT4X2HZBOlF3hGDPLPEfFafmhUYjSpZI
8hkcgcnYeEf0C3ZDCDFBO/4cP5t0NZzgg63dBTQ2uSR7Jg8U+eYsJ09GKNXMExYDN+5pDZiSDIf0
apPgte8rTin2FwmhpEnYzi0FvZDgS2G9V/CnKL9Gub5svc9ikP0V8s2rPI2KoA1gSyz8BSjkOGY5
W/WH6Aomfzftl7Pijgz8bW089+vWGUzE7MBCZJ406RAJ3dCPrwJxhCO0v4n9/7fxYEOBkaHEykxj
7yf14AXjsW3VHxMsnBGtnHPdGyDA2T/OyQ/RvIGHR31P70ZnK6slg5vdl/x50WK5FIE5RLmYphB7
chfLLwseWgS8SD5CsNF7CkTZ1HNEODSAxSFxqYUH5wBhk4tU86J+wWebeA18aSwuk+BuPorMdOK6
VKkKqshcimjkqGzxCTsq2G08OcsvDeiAlIVMg9rUP4LU2oTJ2DTgCBWa6bJscUK6+xGYUeMkh0mW
SN3h9XhRxNMyak3aytLFLtB5VYSu/Dze9HpGNoLdNIrZyxE/BCg3S3xJo5VSq4JOIbCCiHv9HwsQ
XusU+p0Z869iMo4N31B18dYaDBAmn5929CEQrFUn0/hX1pajsq5J0Ovc9kI1tN/GG8UhPq6twbkT
TVuY7Ke5v8J3jR9bFGjdPWy+aUnG6uDOKwV13gTSOt0P/WbwYXkdXbc3wFGFXqKqAa9j9/OhDy0f
csvhB35LGqf1qwKMagKtTGDTMyMtxGfftpyYYXOlLkllz0/ZEN3e9/KPELLo01OSH8VwIa6K0JYb
l6v9Af1oOAHZoKw3jy6Cd4+PIY+pPj1mtEupaQNNfFDk061HwR2/LgTl6NuYxO1/SNpPm04qDoyr
pIC7y5C1go3Lq8Kj5nwkQRDGaQzBD3T87BpdfKfu4T+8fdsNS2ufN92Ue9wFLlWa/lpeeNNrEo9L
1XOwiL9WaLRd+MOoPmOPZQb5m8G45rRNTHS3f+95WcoQQd9pB5dpaRq0n4vPmHAjvnrbzsOUQ5zh
iFWgavx/i5C2Hgjl5ABUCmcyZ/2Zp0qJNmrixCDNGposl3AI0h2EMl7zw3MnRmwJPjKa+h58FAmV
bnZgxFyzpTR4K2dsUflyAR2+ZP+TkFWCf4MYgik2IGj2L2mMB1f4HM9vkp1TmD4XV/ilM1Ut97w1
IC283Ytqk+emqqcdpaFCIuj0VRxb1kVeYJSnrSAKCR9lPs3GmsAGRGXIY818+oRKyQau6kOVa1DY
ll2FdfIRkq0KmL17suT4R27bttAiDtC/fuSrWAuMHSC9aWf6CKSYUsDhMhf4Xd2PwuKNlQWmh7kV
Lt/BgMloomSg3t1iwiGfZfvzKOHMTGoFrZ+tSbvyx4W/YphPr5CiAsMJhYei5Zs/AYcSdBRoP2Hi
4E4ZVaqghu6jLVppFjYhMJH3ULOaGfbZEerpqgmvw/8hbcjSsbv8H0m40C0J1IMleUXwY7GMh3F2
H3baHnrQRPgjaVJND5KgiJ+Prmm0EgQqo0gEGpNNlmUp0zN+S/cbw00r0hsJTfchkLV4nd1hTuhb
a/zBpyoGMzUIQyuQugFJlrAcsBWSW7QRZKS8F54svtSOAziAKlApmVzDuR5rzhEe/1oKsTjgfGpf
cpYQHItPrzpYT1hVlocpo6W3InHgJwBjXOwf9djXptKsT6Dk5eAbMUVcJMizwAwrJUZTB6OWLjta
PBhardflPNHbJ8zd/poRfF1btCKZNIrqg7RtmJ9xue4HqvVITSdHwQMXGJbvNiRVK6vFjol7zdDR
OXKOzTmGd/HYrEnQMZr3SRklID9GNvx3A8XLRJgcQcf+IBqvvirH3JqzTI6CorRpnrC6tNNZV1GX
2AAbsbWk2idU2ZlGxKJCzntTZGEHsLBMNeV5KlMQrUFixVybIyO8v71UFgnjsvLYJWdWDyV+wfso
WHd0NhnoBHMIvDo/J5VeSFeUulKKXYZrO029AHQCo/35jEqhL8X13vsO/PHru/hNMm0Q+X+rtBN/
n70uiiv6LHbCBB2vQCyeblxXABERXRRftOZrUltKnlCPzSj0s3l3vMn3lcj67IVKoqp5CMqbV41J
iha/RFOXoFBwipPGgYbtwnEDjoDEfDu5bXi5JpF9mwnzrRSinlX5+0j9XwpbzduP1OA3pXDjMgq2
/kgthzCN1X1kvXd8krQEZectv+nWsAnvNG4iEcK0Ksd7/pLM8IEtubBGhtPjy+nDNBzGiKjyxYb9
O9dRUhSdt876MOi8Tbac8w69WcZ//dhcshkb5IWEUUVsVGZsM7/arolfI2zUtig4Mjgcap7CQWjN
+TbeiWp3cOnmMgBnxnhybAh/+L51pViTpDBpuSRuN/Kph9qbmJz+1jYGvVEayvxU0uueZ+ef01Gw
WJBNHhnR221lfsbSt6KwY+YhUZ1mULMfphQ0lglpnpIpC5wgLHTG0sv236ee7tCj9WTWSjUNxPP5
2xuW2ttKleKGjWF7kJetDmhzoOhpePV8NgmVdgQPkJjv2x2I9OfIbyJBKjG+6lnMuicZfNo6oE6i
JMb5/4cukmuYV/lRECT+534SvQhEcPX4zQEgnI8bJwQAy2Db4n2tjutf3re84886QnW+4/0v+XLm
QpvEJdpIk5ooBA75CrPJBZ4LpV40fXSAJTq/Mcj+TtuMi1QrryFqF9ACa3jC7wfi3B2nrQQe+3Pz
BouZA0oiwOUaOMXmZ9z++eYKTkgn60uhAHBlX1OnCqoNANsncyYs3L8XnHa0EW4JTCOa3LLPiRkl
e6NaPu+t+NuQ9sowPO3BzCvcFiv6hid+mwV3ZfjrMKrONssRycX0oKjH3cLhWjdd8DKZYCh0W/z7
MxZVVmBBPqXqaqkacD5jf2HCas1kgl2xYbBSTM2stG+WFcnxFt7ooLCqQbZg2X2V0lj/Yoz/wPDz
3aZXnYzmNRjB2n7ni7mkJTlQvuPZN4d1h2h7t1m55cS3zQM9rzov8Sup+k2dN9rdG5KxVLXgjbXt
Nge8wJlCJw2zWo0uvDK3tIPCoYrm6PF8fFSNBEIfFlUb4dUS5uPI8PMwPTLbHBebnnKT2zvbkIfz
sIkczyucrdQQNqu//I3sbZKIHGNI6rcFL+U+84gPsfhS3s7JBUth2eBQ0zV96XFf00pBt+6Ngp7G
swGdJFsodZ5wpuBw8kkPsgaF8I+B8xjBG3bvdfFZRBg5yoi2dv81YcidJNUmjIYt5jcPrTbL6cbN
fzb3VGlOv/CziDfcp43F131Qwyb7H6vOkFIUPd8AQplwewwgTfh5HuMSq964t5FylYgmzvvcEAha
XuODt8q0o2gRJo7/FTXJvQekt6UU7tbW58F3Dmv7iHwUTNk/6sWC3KHcBhmJ1xqdxiUxgj5g1zKS
fYBRxy9k9p2OjsIchvpWXowE9r9yoIwLL/UKsPWNorUZZDgoA01MHy4SaMd+Tt/5TVxv7QmJmUyF
arKRkk63Xl+amW/RV+xTJVbJeEIYbAYJ6MFN781WwdogqJfI3DjPNAAvpNXLpLpxmtSWUAj+Igwo
t8Mtj6DsUJA84hKoyQL+v1bYLqgNMagxapF/j8nZmM1q48onx2tbki/Sf98RUTFypp2sY7bKZ2L1
AgNNOlCr5K3JWHTNLgGMgzic/ubgPoEEW3IUL82W0Yh2dIB/Brid4khxhTmwl8FMyXtfhzq+4nlA
D175v+GCHWWbTVRnMmYIY7A1cZlN0nkVJKoHU/IzNmXyvUuM+dOhC4kVMc+UkDb1A+FmRvoeEyTc
HYT4IR+3G7h/NrzCtI4mT+EGNxGDfRxEglGyuCoBQaxIQUJAKOX17tYtbkc/ZE7o8zzxWtlRUbM7
Nx1wddQK8GRT8ZeGkAIhtaXlkroA8uD8INRevZm0zGMWVaLja1TREK556VITiE0qQcUQyex9Fulw
DAzvA4d84oQKjdsad1OTu2QlpR3+g1f2DCEZNKqNppf/gDEEmelsGyxRO5/Xktmc7BL2Mcfp5hMp
PQt5rfCTzKmsD7LTkGfyGleNmm/jlR/igemdU1EeSKnxzoUIZdxAf2/QLELjh8q6ihPUhAaQ7ySk
FNU8TfARIjoRS6YHl0kquxTGfUXDE5I6tVs0+yqNTgOeOiJ988A5V1frt3ngjN0AhZJr3SeRnD07
UfMKq45PuP8xwNNmDqHdpZi/ZWfe5Ptmn8NrFHCBdAyM/n0va9crrW8tU3OloSWjNxigpQFAXxby
NyCM3w6Pt7aX+Xzks0sErN8xXTzYhiTThE0wQhtdCLMRX6AhBdj5qHIgXReNchBfBZrVBaMZdadP
9ATs0CIERZFMDS82eK4u/hA46vK5kOnMDLsjp3D9TO3U2UDk0XYF5VOFsbVBeKZ+xP+kbVg5LbrK
Z99Js/UJOL3n7frnhl8luieldc7g2d0q/vtQJNfc/iXyaFiRirren6Vx2MOK7jAcp4f0ZvxhXnyy
GSAecuz0HYm4A1Xv4bLKrvg3WnRKxjuL04tZId0/YYCl32PQHGORmVyigJWzyKFbICjMY5/mt4JI
jpdCRa7OtUK/XdBq7GAzupBgx9H1GMeHND5ntvFh48U6z+Yf5UTdPRBas+ilmdsO2lhtNHxLpatm
sKTtLW7VC0QCbg/64sB4Kt6fEUYNrt55xaNnqEJGr7fOBtIlCLx/7dFxQUK696Yz2W1OdSUfEoG/
yeXD9yz1TAS7yYxjdFtdnjyRsK+PK59yyIHYPIVaRnq3+ZL600AyR43SKU0DdMfKZlw+zcT5R2iC
gBkb6I18vvEImojvNzKqnYaedgH4C2GdHQ+rRLCzulCT1Mwr4sM8H4gqRUE+d7QoHI6yUMgtq7Q9
P7Oefmj3XzG60Ws4emnYTepmSNcF654+Ibn9M85GVcG6omhWanE2xB6dMfSX22Hbrj56it44RNH0
7n7HXE/e+gpyJsiZXqso6hMmM7uSeNV6EI3qBAyK0gtZTq4fAfLALX2aIqR8gt0s/Z9XFq7Xn5O5
bzYAeWd3ri7IYf5/WcvAF6FEhgIPh9avlPwflst+DkxWKqqMtsRwfG1UEy9UHt7vzx469ZXlGu+2
29U5HCaXr/KzaDq6rSZkJ038RU+x5TVODt5YdUAGf6/kkmxO74taIEFw8hUi/SZ2YePllgePRvWi
1kx5c05ga/E2UlvZXF3p0Qbx37f+T+/462LLTuycV4KSsJjAY0vlwwZ4b+4VE+Pftf6p2smHmNuB
pwz1i4h5D3BYQDItVHgVa+0rMSF7h8M/4yY25AlTGT8yOkHjh3NAjtYqOn4EjuISFDV4EAcPMmOE
iKE5FWjM0s3N7dINXWTNb1pR+E6aNPi4K5RCgQXTRWyNGEPRpXouucTk29VsXdZLs3iw7XKirIwK
MU197AgP4QrXChjd/s6hdpIYZMbHAbyOMIyOvFYXh4gvBzhXm8+FyZd3RrMP1rrGWh6q6Qj5w0tu
C+7xZe+YZmDVY86bwviae98XYZr72SMsRK7/ZHKMVTfL5gq3tDsse1QQSDwqHwhjXqw/4+4Cdvf8
3zlHgSBRTM1xpU2tACVERXv26GMNA7M8jDjKgl4CWN8lv0geajR+rSF/Gz9hMPl8Ai85CqSwU1JK
V88iwllIxtBRwqJqdBTuA8iGke+XWMjKji6JmxwUXveu6oBJeK4CCG56ZKBHdA6T6A+md6E3XRjw
E4mL4pKjkq+WosQoTSRAdh3n5mdkdp8UCneAQeN+u71eBA7CLDPwS/HzyEx6npBa9R5yEkvFkFTr
YsObBFnHJyEROLXUz+Yf6Nf9ECltDrYdhhzuNsfvvov8Jl80SulUyJRWFXX5gkwMT18qr2hNXQXl
VUQjBPWV2y8/tmnb4TkGVAGunMHHq4e6mNIfrUXLHoNetut9bHEcsl/1nN5BqswPzrqIz7RKq9j/
x2QKjXZNZqqlnQLvNUI0DmEayAERfTtw+3tmilOs5xR+qQqL57N79YNW2XGFyMRMMoQM/eeQSiUY
wYzVuLxmL+kCOqSVS+LjYH1FZfnK/Dq+ekMquDQNCTYHSb3hEO4EfSOtK6OvGYAfagaoalwKFXF0
NS64IKaKI1XzfqJQHKgFiL3lEFf6G6ykk8iTHeIAKmU8fhOPvt5Yexq9y1fW5Phw/KB7t+dKEy/N
rIVJMUwnhBHkVGuWcG30WXbkmXpxRU5vDMw1iSjmWJ8fCd6xp3FSg1D60/P/0yXTNiN+W/ou9u9K
6Up67uNW1N3cIoUXXm8NPw0x02FqlEG6eFO00G/ucj/BmMvw7m8rq6c5102TWtQKDd7l4E6mmKid
xj7kZaaUIJuCBmeHdM9dwu/JEoc/Wdzo6lbdn8P5KzRlyYELuSUCKV+IFw5pjaarwPZ7EACJEQtC
HAUXpin2WpZXjOFZxFL9o89yIvgiAK/6zNDw9UdqSBpJs3yUvP9bIdaxRWrPd22C02kEX2Nwtav8
J2Wylzin556cye/pvC6SNDO9k369ibju9BOuummjXCAMoUGk4dCgVEHIlAHZaXe9IWbXN+UTY0xf
JZHHs0V/VOcCUy2KuxLhFTOYyCk1tKyDf8VbVu8kq26zEFAm/wXyLt83iFcfrlz2Wa2XIvWAt9od
a5PWkUo8cGBQyV3mjLUyqlr9N76JhE/frz82Z82i3o8BCXuidrINsgx7nvj+Kvaq8xronlhbNePS
AkgswgJOWB9w88TJJGdUyy7s2JIe8ou6jpWQiQw1uDOyi4PotRngkMPFjp0WdWLX3YY8mT5PKwxZ
H/CJmikY9XLWaN/naZeHefJxkdlsdmkzImoqu1PccYtDuxZ8eDticEXy7126LtNz2z32lz7qr9iI
xjatNdH8iE7ozdSDhJeQlruDajdBWkt2eYzSkGnnPFTyd8KdyIeo6GE81pJr2TIItUC7cwYpboYZ
eCbS5sh1/+k29CMIyETSqzLxHR1T8BbcqqVuCwb7oHP+YIGjBgfAuuF3X+Rtt4c7gCiAr7clGKhe
U7B9ZiO8mvxHTfS66E1lADFuZD1576G36eimbG4C+tSdANbNf0luBRySUJwRbV7tzDc/cXxk7cZ7
hc3MH7JKI5NFw7XvrEGhFyV93zWUqvWtq+IVwcHZhxwh0n4hNV5ydnpQRbAKRjTQg+f+uxARJIPp
JhdwIFp9lUOMh3hK4Tg9weQVLjhkffplgKkCTqf7wd7oYOfjCdmEz3Wj2XvkRMcRq48WZm1F+I78
eX6qfEB00Hqf2uSHzFwWnPCYXvSEJts3baf+1wBySZX9D/RUk4SMyXsEbinhYAtXNB668t/IpfYx
p/WVbao9dYZ8W2gqwfSPGLhY/jdhr5UtO5vuV4qhCcrZOhOvC8YGK26SUEp588BM+pBltSkWcHJf
GbUIh7jK6R3glJg7JNkULVPhQAFjKFzBUfcR+3zu3b2n85xPLQ4wOYhRL8P8/vejXXo/Ii3eUU9K
Ce6gK4s4iBO0xRzhR2igCVvUKNKiWqToviTgMqE1bWLdHWINi1DnC/6QRB+Bduc/GLLuzYiUN+67
VsQ7hoTtNkTGsnTPld9JLKAyBqzHLMAp+j2H+73YJEx51rLRByzpgOuvc726Oje/u9T/ESArMLnR
Dhb24TCSSlJ8oGF1CEB+NMB5peQAZVCLrdy9+ny3A4jkO9UpI17aSREPTOqCRhKYYysI/+K6rcjG
EHOvasbPdb2e65Ix32j0WtrrH44NHIA8JiEbAX5XpT9UaGZ7w3XPt8dOScj5OiIT6iuFDCyafvdc
UAsAecJi4VsGKZsAV7kLQIUR0Y/7eBzL+A4+wZRaus2rAetq8RAeTTPihIAMOWoQAz8jvT1C1SAH
1FDpZvxq+QzTvZf+9g61zI/1cEFfmOTjJEEY+mKdpbLQ60sYLIudlflenjEgK00MtiSagg8KEsYi
8ugtLXA9vFjGnJ0wJMRsWUekEWmXQ1CHKuvWhUhBPFWcdfx+fNZKRMhGC7cexf0w3MlQEDIFRi2L
PIghO3X6GF1sNdgzXZ0sHFGsGSX0HvapyIkDuix3yK3jBWlTT2K9ZmcFQjLfFCuysLjXYHAghgOd
Ov2yCNvOMfzz5SyTQQRUX0T3dESr5ueUDfSUK6SHYiD73sJx5s0IlP609tDAHjcsTK9wHD7DrklG
ZV23dswrGHSCgIRIQXRWGLuaTWMjHGEn1uQjvKC6N7cq0eiDTk/dEzIfQnNauMTAN1SYpubDxFD0
Lkv28m3e8b5KzIhjhegCiM9+64P93iEzg+vtzwRGW5NEuDv63xyqWTnxeBFgb9hekMoanjBGZs1e
htkxgyJ/coqBaZ0AMxlrbEC6IgeEnIzkZbw8XpMmwIFqkPnN9NmsO6Dh5RcB9gDvJW7g3Exi65i6
QVvfTHehOQTRRNWzQboeIcOBduKO2LpibRJ6WgG41mQK/wq8mSUyysE3Xkpr1RObkrxeLDHaNLzT
B4Cbj2KLIHvuIlDESyCJlLRIdR0B6rCT9XxQoAdwbY+/jdJmZHKiKViwGd5m8VmuTbglfVSoWaVp
Qur3T80H4WS1dQvHfdpDEiAScCRozgdijIuSCsPmzLRoqUXDQ50VwMKWA9BKGW7YI5B7WUflNQCW
El1mhJJWFiJjIt/nXenjCBpfy3xwp3HtVqs52e7lIu7+cx0cu2eLR6J7U4BpUtITZwMQyFZ6b8aw
mTkxMToRB1knUgRdUeJ1u11hXN3tWXcrg5j0Q4mOV8yWn9W3vp6SYCrvsvDp50qChO17pg63+mGe
O/dkfOCiKLTBrbPLIqT04XFfAhoAaVJrtmD+zW6fEdOS6MCPri+E04iUMLx9KY7+zm/UEjzpvoBw
4dlV6hZh0xjx7L/FFjnhD+qnQy6OhPilQwetxWmu4yl+dpFJ6a4gGTLaOnhSWgba8/4/Y/FxQ/Br
NyYlTYnoF4NqKDtnDXvqamD2o23tPa5lduFsnBE9Fus8wiYFlBuI1/sNl+RoBNK5MF0O2ScGTV/0
lPlctpmfslkJBMnkQAO0CpCvoshd0U342kH772zQLcWzZo4kuTcYtUC/rDmN3051aldOyd2xKbzm
Etw8LS9Xj9W/eA7vQEdtE3nHWbAfELg4mYdtBpREvtS7eroJCVpjrtXkLWPTh7j4TZUHkSyBU3mV
E9Pudlx3PUWygvp3f3x7AcMQpLotJnH7bEFd9wXphbz8YqlRyoLMkP2e0N3UFTq1G6bjDUq/4xRl
m4A2dlGryeuQ1khHO0UiEc5GVGBIU/B+xGgWqTwbGQeqTo18kzhRdbZ2xRiqPmetbogZdidDQ6Pt
PoO3SOJEB03/aOcXLeubxhGLB3F+a6GiCP0ubL/ldDxoElFXBSZdxNty9DvRGCEDoFE4C6K5qqdn
wNF6Ugf3ggry009UqNsZ87zw8cHDNiPyZNOZg9XMnJE/hRrOPERYWFRtugPGat2LkGqn2i/fHVgu
zNmUZaOoq8X548j/YvseIr7T9R5LGrD2CdR6muoYn5hgOEcEdEwoIKRtf/KY3wRRy09NKVRvPVei
byKXiMHQbABdLOrpZSjyJOywbhtYeULJpmgm8k+wUDQxblfmTK2nyXAkhaC+E1TyShyULQZEnGy0
waPkZQN+N5sUlG4oXi/YewXq6IgxWY5kYwDDKxkmJKlM8gy6xjXSLIjbLBMWCl5XJXusthX6tfbt
IZre4DNsd/OTS2l0NiuaYV6eEb9UOmCgqtHHaz9l9tzyCCKBG/Fi9+mGoDcKjhFFzooDYChKXf2h
qXkhGC1HwEic51MHb1dDaXFdrGbbwBnD8ZN7xcMWbXsOupCET+2DCKRbTQ+AC/5dEN+qk5wYeQvz
XTzYMrFe9oQzHsQWeUdCHTIeCF6XTwtFG50VAPHxAbVgBkX98JImWoI3WLWSo9KoL5KcvLKxohYL
4jPvZsjjlMRyrTAKQth3laLpqQUmaNhYzyUpjyJa0n5MK1DYJ4JkB8w7Hu7Cv+KWdaXjtgsLwm5T
0fHEuOnvxLhWfFxskKm+nikGS45X8g0rCVbMvXHo2py73mYRUR3OQpxu72dXeOf0LogWxc2jNsAD
wT4TZOOf8VilKGVJUmlbD3BCtmcubcktPDVoY1We+IhLavKeDYHHYqg3dIsUujz1UgBijkCc6V7e
siVerYSR7JhjAaSKo7pZ8kYgS4jspXQO3+6R467D2JOOJjS7aF0r6f3X38/K7GvsHZgeQ9cI1TKD
v4WsT3YrCyFbI8oAuG6KPDNRTB+w6bhN6dp4/k185HqKi5P+8BCB1dWKFp00ATjCHUObhGhCJz4m
wz4tbHOR1Dh0JaZ7chDwxDsEcDlpYOePfccUNe2ADpXSlnyA+NTnoYxwn/dHKBUP5Vbi/+enYHk7
hjqSTeVLn6muR+/VcNSFQzwbDmdv6QDeXQEKS+8wrVjrGsDx8M/vMzFxzpTl5oHXo05PccnvIXwe
DlovfIfMwKWuJ5ab5qlqKhktuPnEpy8K3L1Pyu5QilhxITfYNqzyVvMMVLIKS58j0ZjqrKc7M34M
Xsb/ODGgb4qkhw7x0c6KysaKNMmxkpZ1f6v+1y5PC1i/mq1PbXQJhY63JSmrAN+YUxozvWBPEZ6K
fFvYboXKjV4t40JKl2v23xQtdbO6heY9DBt/VZ+f3glmw/+QxZgb2ribzUSuEo/IRr/RMS4e+ig1
danUYrJXtzRQffDDavorUbqsk95uPvHWzbkodcIu8qR/v6RdCrZp533HIPzA02HonbrWwq9JQZxA
Nnv6pQof75ShyRSuYwlSTYZPE/BZXGY0x+KitDNOeWCPfgSOd0LZWnbwsL8mgiD8DybyxGS8zgh0
TJ26xELEyRgZ63xVz5XgRWhGSsj2k2NsL9vnS9UBLPWqW+qKiQrgX7HvaFk2XDsaEIEFCQhsFsjY
CkVzeduqbmLAtzAW4vYpbQIISuut0wEu/lBoV8sNm8yZcX06XnH5Csn1a/6mX+nTm9f4nQ7bpdlC
UgUp+ob+2VMum7tqpdRkHJR+72VyhueXeha+jG4xfaxm8+84zLNCJ/mkeorZdBeM58Iihy0ouRn8
3zfKWxqw0bpdRcHRUJ7T6MGYeLgstQ5mGIhnw9BqUEjNYkCKzHZUswpIoboFGZz4kXkrfhwUt9rQ
5mEheo1RJWE65JJopJmrouyvLbfLFni2qqLIT5Bd4Xd3KNvmG3oLKTFphC5A4E9jInx5H8HbUCk/
AubFEQmOEwT1kL0Gmxcnfd8z7t94ETScfBNtcz1TUwvX+w7T+iRF3gfxJaGgPURVH1UkroJc5DTv
LFTn0fU0FawnhopDRx0lAkkh8wH/3jI6xhC6RJW2BFIGWxRfMQJCPh3G10witUUo1J2x0DLllxHj
+w6Y1ZvsA32f9B8KGFjGACdMCYj8nC3w+DC2kY7PNwcyiCJMWph2l7qKiQhtU7mnQkQXfc2bIfJE
LnN8X2YnOXeyEjh5NjQVvNtlCQl6/3O6zfvxT+Y3IdMKaR9400nZmTovCVV3PPFhQpNazE5wapCk
HjHRzRVPds+uL/lXq/l3wE5T4SIKx6MvtTPdnk6qrNqS/niOJLl9Q7eXNC7rN+wqkJ2JGlTpHtoc
th13rTuxwR7nVLPoT6rv9m5NjrDMKt2Jj70hK+/Mp3H+/g9opYcz58OTkj4tC5jtGtDQ6evKjvnM
scpnaJkROg/On5RVD94JCrvvVmLWjYH0QI1vkZIqKvbcOYAEhHCSPTltf2T/AZ3WY+suPaKlw0FC
VIVpgpRE4/JW+KeIvM19m7q+3I/tYGpHOKbfcsNtukkSEMGeNFE8gfAmlVdv+f1muR7wzNeNtmzw
YjYLRU3FJKcOJAFJ8fdkhC8R1uFcDKh58Y/iK3C08A6s2mh5nI0pF5OCXjHwDmBsBXT2ut2Lc/hE
d2Ck2djAu0tV0WsUHymYM8/IogY5aDVlStWG2e5gEhkD1f83DO8chsXJNfWhT7NaICvHUSYLWzWC
aPvnguzw6mUZqlsimjcZjwWQ4iJgmHL+u39GdJxuEEldjrD5x0rbFGCLgaGvSpWb+3xIFtyDw/7j
bNdI2ocIWf4f+05cxZQR8TUvSVY6+BuE2Vhs2x8UYmoOP2ycVKJ8O6SqR9tXuIJzDuKEZro+QUYs
s80MkloWgsZS86BtoPPRtCV6llub5OIr+MuD+K5RSklT/KfnQgCG88bq8v+gUKWfyvRw7DlIfPFk
xvQEo4v1QiF+VBfhWUoPovAIVSISOJ8e2AcVLc3HjzJGgll0vi+DhnGXn9bC+vFyj4APOnGIOjX4
fhx8plmRu4pLxQPInyxiHxuLtaWd0jIipETdHm1EiVpPQ2u+PelC2388ddyQdDDceMpDhjJYqcC8
R9pIgmpsbt93rIj2YhrleliVsjXqAnCLsyHpwxuaVlhYbsEaHa6lukKDXvkhVU6I9zWmCbrJ3DNz
b9ElQTYy24V0I6wbmh9Ae0zDr+qJvGXINyUoI3YnNhxCl+J6tM/QSplYpHhurdyf9ZS3xaWCLkwJ
LcBSAHjDCCHUUvrrfdEo6BU4caEBuQA7f+Ki0LZgNWhKh3YbZbPaBupVAf1ZySwZONUR4KaGeM0M
vMwinCz/ARCPHX2T6b/vNZBKx6kiTSJCeC3u4qRK45XKFAZsKLyvf/6vAYNgQSJbrmpCrilSep5a
RWcu14Xu0hkaV7FX/JbreJRVADCA4IQVmopkqqGAdqfc+kLmCdUFy72msqpjkYDs6adM/vqtxl7W
n/emsb61KMzSMF8o8hPZTbTkNIbS9rky8DT1+S7QpSrYlVg1nPIS6PdBmGitDkknK23F72SC+Wfc
6rJyG1xBh7eCajgx9M0GUiU3AycvE8T8Fo/EqJVamtU9MNG5fKEY5hBQQuAa7mO/HOdnHwn9C1e+
64AG+WZhco2+pcTFPeBGqR0cwrd7ql19OMz/sr1R/bOSt1MihhzaZqAW3lZmf+aeLj+wmisZ9ljU
1IrRq/V4wG1XL+HKa3DjIWfg6OUQpELzBqRDy1Z9ComgeSVMLB+dFl8tSlIV3nhytOhNr1KyI4WO
5rfH62Qq8f557Y7MY+mDbFqza7IxdCKOjBhvJsuPnsWfmBqmGZGYQiAVKQXTSywZellDJUNK0sf9
fuYw1GYKuGUcFMzW0m5e2IM7gzY19jJukn/srblhRQ/+YnIDjsxFdWBlw//g5S4jo7OfKIxK4yHn
3Ql3lSsQgqAFUHAykC/9EHL5OGi4dblfwP/lv5YheTY/pdlT6f0w8/VP41B4b0nDcb706AE9LYI8
WkD43J/f/GSKBkdv1CxAzVv3UEhJ1CCbnRo5UFSjOYJTFvQB1sovIgiY43P9LDHvd9Jc3f/zbHw2
bs6lXjn6Lj66AqO69hFrO5JJLflc7FudO/Ko4wT9dEa4fpgWaT7bP1/Jr1ZPUi5y8XBxE6T7t2NP
1nQZML41SboOt9//Zk5gRq2oDsafGYwUpUasMN1liLYqoX9bxf0zcQztxVKL9RZIA8aydunFZQBL
mLiK7UDKKv+nEgwB0Xb6uTucVMg9CbdaFTHD2BkKrlRi2XT5aIBoDBLJzsMq0TbhQXHvTCXJ6n0J
pb/G0Gxq/8ETME5TJw2qjrwXWr1ATWmKJIaKCEZ6JOgf0GFEtZJHOyVE7Ly153J0t5vBN4/gR5vA
7pn/EEh5wTzINtoxtysao2hYoNnOSOwztGn5VajacGsBMTMsDFfaN56bmjzMD5HzcopeX/aYcTGR
mMbrKiZsEcjkIZlcVEgGsdAq+JWIgmVpiPG+Eu6sEcOc6yWk7vLttD2qH9xFqIoXmAijnkXo5OL+
NSkU0HSHNFVgjcSM/uaeVhO4SSuKP/jmQQqjA+3ivoLE5n6rePcZ+GaTPpbx/n0GG9KGcLWo7UsO
nQLihWEXJGIa5ZHpYMCp7Lb1SdgA2OXNu/FvDqSfnWsmTVxY/DhB3O8DQaGY+ODpLVpyqhLrL9cH
iCMYsWFvsaK8wIDnfBX6W8DJdOeHuRscROSdpPQLfoNqZfBwtgcvCecIZmCyo+kD3KIw/pDRS3/B
cVxHi6cBeP68QLZOu14qEFOiSwa1v/3u1+GlcmryK3wkRS6VGzBettVqduVp79GFVmWqnWyi8s8f
zs6ZaGe5HOIUwGiEKcgyx3fMzSDaE2NK8hZ2pfkbyoq0fZTUHM4jqG6dvDVT1fGDQmPz7775xc2i
UC6bz4vdk7wo30p67ibjg8g1cauc3O1Pq4l/JgyVAVZHA4Hx+BrpRZUC7JtgIxep/OoRhnUSOp1x
o5/AmSj0X0QZLKwxsEfyKQWz0mde5htQxhl10pCzbTF69FTTSytBO+kbIVyJ/pcYYz0viotuRcH4
qmYrp0vHrsN1aI4lAGRlfEmjb1eNkYPPRcOLqPndxqoYXGt7h9/M2NCKEvzwxnVYNFdNp5hmxv7o
Iphr/y/r0KY2oDpPq52VlzBzo7R4EQi57XuPk7wdWhkjiGoXSTrbwUeSa3cB0cJIFpfr26C6k7y3
p1BYt5BlKChPTgwNZu9RDYoFRMuvkaxD+aVDj6NGMHBZGQ+zaY06MKmvX3ne/zbxFvSOjsiPms7O
hSucS0M0pYmKn32QGgMJMMaCz+6yh8e6v3nkJZtVqA83sUP9NCNXCkP/jSgHRvVMOlCkNd41PCu0
fHkIOplieidq6BdtU+nZRYPbIS0jbcbeuA+T4LbAD+xPR5EZl4FAFvG3C5evX5ifCuVAFHgZlFWP
WM9anf5fDL8uXe/k/n8y82JMY5T039J0iTLWZMimT3PgQNtsNdDF0mH97EuyPNRqEN4tYK81oU/P
aKWGUeul1qMT0yX+5Ia7KfYULf+aEl6UxudZznrkl28cPteGpKLa16qLO65rcyUvJo5wZZKvDkMU
0hzcc+g91lRDXQWhphhtfhM0ATsN+KdGzlTNBccnBBpqSHDajv2+z2XX4+NFA+k2yXgpFsk49v0u
F5V1vCkbpy5OumcgOAfPdZybjUifAH1dB7tkH6FMuDHmLvmkAslm1QZf4m1+/7tgepFW985jAr9g
D0ZiVaid8NVeYNpy9e5xHdBKj+qCMZWMtzVtGi/kp6SVgLG81LmQ1JgxhNR7JixVxcfPNsWhYg1n
IvvYk79HIdYn5AhZ5Giln8tA1TqLXF/zHIMQt6FpgvCydx4jGfavQEGeYk6noDzPe9jJzkSHnD4F
Fs2dDZCuHK/O332kpXXMN8NEWAiTez39iz1O8zrabz2os+hwhISW+cpNCpi4pLIWFqATHUIAEv+F
keNog9jmmOVVPfR044H0tgrwT6OGrb6OEj73C2SY00LTBpgLXhpyJ5VPFFd5Hv4h1Y3ByVraD4D0
5VhNcmz4To7QmcMQhC3im4s10ZUl+HJU8fiCiX62Iy92mHOWmeW/GFJRStvZ7yRYB771vfk5EjXe
715EIk4f4QD88EXDp8LYRzB6eYoJkjxqcBcskaz6RRG49aSaKsadRMowljRcqUiXGNMDjifJUqT7
tomofNPCEXndqsALEs/9yKLHsWUOaToJWsFQxDjXmNT7QncYXBkGT5oTRcyjbA54VrCOMNKWl+6h
MtY0FLQJhRNPZ/x8C5godvUNMMSw7BXFiALfxUgn/NaAM6taunYM2VSbusMePBfb5EucwDGfMZfC
lJB779JQrsQon1be+ogEHZLlaJZTzSmH7dIvu9MK71ekvriiIjj5mIpDN7ggYtSGxeQQvLRPpyFv
gfo0EYgaICSD4rTqZJs2/2VxNe6Ud6msrNRIERfCEd4BE9USRXXJeVEIThK8/mz7SmBj9/zkkuW4
9q14a8fFpFgvc759sn7CMdVC1KsaJMuQKZWLGnVUAA+Mb6tRLU/G/+yruL8Ch1Xy3HHD2PmkipQU
Um5UkOxYqte7Th/AdIelMlucqSmbymoCl4VHo/a5gnQ7u+DVGooJm88QXP5bb5fbs3wqZ4IhBD16
ngbCwShR6FnzqZJLW+1UTBYUNz/wsrZKYK4y5E67enqf+jw+gyzTHiXZAz+Hz7TXbFmA6Dnd953k
1G0QpXuTvYEkRMhedBcR54yUpaxCnl60KqbeRo7di52/3wWvBIvXDe3NFP7I1BLSt72pypnsZvmR
HDSGWx5lvpbEwkj8oEIcVq5NxooUMP2KYGCAD0bnTtGxBTY+mhOCbdIbbvcmvCdaD6na2vWkJiyF
ohj9RTvu4W8ZHldLezLXkrzW8/8jEqsperNjDe8r2qvV5usR+OQrnivHH789RPI/4F8rAX1GEGZX
r2dQnjKPE5A/hjwo4v85VbJVVisvKtphnSU3fA+AxPUYbApSShrkAyaMEhRcg16IxvtwG+G/FduN
7iCOTElKYtFeCCoxi3jaE/+GUqb0QyuFHqfX5Om2T6EXAdh84IcQHPjLxdRhLAjgrGyt4zCS9wy/
fMHNHarnol0S2ksvy6/3VaffJoIzuBUWagsJdPD8i1Ndhnh16i6GIc1l0PGBKpku1YyI6Mk/PXKP
ISy2d46lEa/Ksw+IJgwxgx+NfFe2kiz6c7iea9I7cD7ty0xdO7vLNM+ZzsCz2f/Ly5iHlRp7gGXM
+ry/DiEZjwuKv5Obe/BTcGBKg8SOJ/4fkhXX7WzOA4v+UJx9AtextGPWgmokCkqt939K9BQrp7Rr
lmutESqkLlw+JGOs+RrgjgmFn30bqgAQ9MWay9uUeTrK92MQFR8xw74AOdVUmUrg4F/qZMFI60Zr
gzub4b2Tfaz6xZmZsZSnZ7sM+19qxaEVVu/7NlN67qSKqYzfjKiFYt5/fJgKwcf1q/lsNvS36WWF
S0vghel+A59WTO6YCRkTt038MTrZK55b5g7HEC3a7DEVY4hVmqqoBXt4Kpcs4KAxzg0Cqnwh5AvI
g7eBICdmeoKE74JlGt84VnqRmbLcIVoTpsZBZjLDH1t5sd2TxWXPk4aNf02MLPwhE9eHUxtW+Ucp
TKaQJNoM2RVgLkNv8ijlTQtlygbpyq6IG4CzZSzntn81Ix1nAqPPzLLEDzciGicQV5O8Cl0nMPC1
OYaGBg2l9BVtUpBNjhZB7QTXEWyQeXuBV/ncCeSBA9sTbuTglCmMu5IhB7xl4X52WQRO186Jk1gq
sxZKqX3cHmxrYJBZw2MFsO/jvQqT3Dj5WWgPG6eKZ9xW0AqFwHo+N0tiARZQZklKQASadLYUpl//
edEgka6xHpUdleb0H/gYeMRINJpwIxGOeQnXmxfgiBKiZkPIHEIzDUH7z0jtPhSRRTLuLkwk7sX4
svNlzca1E1pgQMW0n5LtZAzz6Vn5Tf+9IkThrvuf7ZeERHT5OQwf520mbCPRBIsl01w1dPd3mdn4
56AOo6ABFHvRKQRog70216eNGeHGTrsc6wrft8bpwUlGp9mTDMGtS6gIfltrAukCD5b2Lxb7dW1k
l5cDUe4vmeR5v/jRpP2G+dz+1D58onnXWAFyImaIBsJiiNfmE9lWjqdESusrv+obC8BkDG0BOvzz
uksPxFq3R/jSZkHcORAz4QZu7D0LW1EIWEeN3jmmZhkq+PH0k2Cng+FVSdn+R9Hw0NTXYqD2WOJm
lItsrlBKKyPFC42lBBDiArDZLUlaatvIqL31VoWM/exFwdnNqj0xpNhovrvhNUJcUHC0RGRYxSD4
GQvjT6lHcThef1LGPz05gIWW9V5Fcko2dMyTJwF7gMJ1mIQ7pSIC/jj4Zxdpgl3IkGquj9XoYaFJ
UwciRxTDfRL3NHcpRhnDfgyO91L5n5fuBWLglaRYyKvIaFa2Ij4dvKSJG6obi/3N7rPyj9qIyJv5
1z7Xzr/fHa/Rph4oaPuVGQ8RmGhnVnqhjJtzsU04thkhf8MqLsf2v9Ir8f7agMIR57B119c41GO5
XEq9vdKGQky/MvGdiJKWTn/bMHCiecq0466qBjuZmGSf9ygmGgRn61M+DxKK5dpAyXbO3dwErN3L
aIoQqGJulv3D/yptm3oxiQQZyNxTCPOUYOUix3TMQR+os0TTVnOe7uy0R2y10JaxT+fV8lTrQ7gA
wvUKlt6PMn8bpS3yjrOn11XFDMy22OsgE0PZjskt6ws4GzJXb9IEZMBgAEiD8C8OnFzhCPxg2VSV
/g90w1W1aHcvv2rK0FtVh1VOXacH5ojfNRTNxWJ4pchiVER+5om47KfFtJrLdyYGwVmtlrcVz1iC
R/6ysBMXT4k8rchQEWncUQ4qZ71YyHp8s8+8ltTzgDdhkWDt+7h0UjQbTkayxSCQMhxdBn4HD3Q6
i0o0s3NyzYRCRL/wDqmzIbi3TJTnsn4dJtIAbG34VPJI7uUKt/FQZV0tIrSxQsfS7psxcUXbhp09
gT6CsnJZUkuG5ZN0FNN8oY1J1zRCeVZvGJNRwcqOVb7INrlnRqaZBKTnN3Envsq8/lVehdGlmeVa
vJPNmBL9HTM2yDuuJMFWkNMGYEviKRBkQH+IxZbAUg1f0+2KkilsWesye5l2jFYsd9cE/unszTaX
qjb3Dj4/DhObQeYotgUbnRsZm6TLszCABZxBhXqhFqVVdpQBX/9u6J+4TCp4PLk7pCqG4PfrX66v
oT/Z6fcO48ZJvQHnO5SdB+F4uVMwgIIC8lRRpz9Cek/H4DJGdp56erGGUEU1bmqMiUnyAakriufr
DQW4QP2MsCB5kFkcgypG7V1Hrf/zMp4y4mfRNjcdbbUYab4/G8pxMPRQRjFo1JfK1gzBdT9hdGf5
sNE3img0cZALCnCtqDkMibq427X0PFZ55bTH0WMnjQTx3ZwZyArOXS9jodkF/c8eMZafPyXz06oB
CMVR2gDBZIL1Q9K7WhOBVic2Ap3F3Mce0ZJiphX0BknNWbBi+Zptw/+gfQvChm6gdNClvvIkHkex
QNLsI2fBTuU332tI/Oj2Bw9RAnubEMO0FS4oLs2u+3bhwTkR4ZWnSbma5dUibsoHNAAIHIz1cURt
qdQq//kzfwolcoFyZfMh1Vnh85VmsArgxofegU1MkVcY1saLEX7sqNVjjKotDUQURs1Ths+LZMxq
C6+0qM0uMZlpWLMmd5bCYy7LicEH4DVJxTTXOrmMrGui1yqzk6Jg8vPtLtRX2h4pEHKZ9vzG7y6c
8uppjhgvWp4rxNgyrjPz5TEwOch85iDotkfW/s3aG9049zjEC1M6Yl50ODJ0a3U3GPlIVmKh+E06
SvU/RbcoVYIJO2JxSsFvknYV7b7Wo+EFu38zYC4BEQNyGLx10/SkeHXL+S0bxQcgc0JUVa/w7+BS
lDVYvcT1+Kw7EJlorbYwH4Z6yJDKAkwIgWFeG8Qa9WH+h7VEMwgUcQ9xHNPrrVarRHLhWV2dA3KL
oos/28o7bk/mS7Ecl6nXsxPDEPpertKgzThL7F6HVO13HyAR+EoYfacjdcxI+uTcIEwfz5h/fS+S
EI9HCTvwrJih7r+kQc0MwZZCgamSnKBxDozsndh/lAwbEIPUZr7v2ygFzmnYh2BK32ZaYGsvdLWe
8SUJR86ubO9HkGApLiowysTQ0aL7ciPyuHzhCQ3msYUOXbY61EVEv9wo6diTL8vhbkp9Vuh6rocD
dE9/+oYgxLer5kgUc4YkdD8irl4y3b/+eQYYltjnFcuH7Yg5FRuSJoC9JvyPWRt7ihYS5iLN/eGS
2AvoI+lCOkOCkfpZUWUv3BDaJ1xSh2spEl0IItkUL85l9o0tweCUmC+fE0N2mU0WGaCDWhDsp+WZ
d64/r/+peNFIbCdgTet61k3Ln1RekASLWMfJ+RKjDrShfAduDoLSR0C0DEELT2wxx7a0CCOsNAp4
rySEm2OtlLNZvaegv6RSjs/IFKi1S5bdlb3rb1I9DmqdkqhkGwqoIclwBzm31QHDFptcXcKwvtmu
jhJkQ0RzhIHBg4gHDejS4nO2TuHm7B6ZsDWoD5/DvOnizB/OB0i71sZJVvVtouJunwVeNr9/PDTf
1TbauVmbuo88eQlD2iypwmpavMATGxHuITcT7K0g7zWju0r3ZBs/CZE/iEhdaDSBAQphgotRTrGc
5w+MFBnuqgYm5CjsS4HUDwT/uscvmgMTLxfa1M/q8xtjsXe44UMuUz/YXTPAoGZd0aWMKVzlUtz9
rPJTi/MNjktneBFnjzewxm/pS5MyLOHXj5I3Bg7b+u9J0UYE8nYl5J/n9NeLKvB3DeVwDZ2+lBXU
lPdYsJwj9VRx9lXKDA/qcjExwkJ3BT1ImhyxTd/sjjwYLf3jGj3SbMztMMDXJn05kEvXv6mbqs/T
RluEBUdIjV4jW4VFdS0RrVljX59mo4la09ZLi87rqb42IHlV7Oqkw+KU7MVxNW2KfVevZvaiHS9x
XPd8VLhyvALRgyDysZqa8/Kz275/ip1bNYmw7PW5+8cBLjDyOOMs0nHneA7aCBGWYpiuUxTLIccP
q4N30sOyz2TjpwebN49bwpv2O+AuG1DsqRgZwdd2ba8vqAvnB2Z6mVrw99WF8DioTGktK/o3q7yJ
JtoLAtehF+4yIvfsRFMmyGP/zZy+fNQqokdE6yD1jbrgvuw6bmiJ7Xq468xhq/8dJWTEvYYX2Hkc
CvyD3tX5r3XM+8QZwi8owgpv7N2ctzC9Q4v8fx5S3PVMeC72cDotVLyF6volpARu0h32TUaf0wYL
fsz3grtZKMfR7jPt0oOeRk6WsLXP8Frsjrsm5XX7f6W6K58bGplWReDR4NQLrcGC1Fk4Xf5rF+rp
kSyUQGnJR4ib/fFUG2E0JXEhkvn3SXKCTQiWd01Sk8dT99rEWa2I6JF0vTX0a7hLwdX1tvU3dFDn
OP+uoxDk/8Y+7HVyJ135U3eqk5FNxBLsJNjdhl2+kpVGc4zTPYUpJsApRBF/gF9WMmOAeZwdzhuO
cJciL0Yw7ZBgvBwcVervhlYSRjpj4DW5/Lm1vKs2jg1QRaFKOf5K5tPRJTk8NXWE4+DXTWJZeCkd
R4ncc0mmV41Nw5djtwp0bRLqNshPlojTJ/y0fKQxDtVIZgMIKzanN/BIZ5xiXZgY2OAAJV/BsJsX
VPY+pKRPRY0pz3EuIi/bmtFooJO9p3Eu6XZE3UYDU1FNcijQKUnvNe8M/iMZVLEeCxGM3qMz1GMq
WAJz90qCfebc6QndfxO7cKI1rDu54wXlOz8824oc7YwEREP7NkEFcVjaVtpvahCTXTXVHhp+E/Xi
M93vTFPloG0w8260IhzoQvD1VQKTOMfQ7VO84reUMohvznt/6+EetMM2vp94pN3cnXTg+KZlah0G
kicnLDA1iuvBu1OkTtp8YOPX/ot+T4/T7fRBNS3yNBTqUNWTzUe2TwdHFlYgvd7GCwJ5zqD09AgA
EcYARLSZF97KjykOVXQ8vmQaLlX2amh4lS2FGw3Yw2KsWeHbZLS2/U4wzBm3bIImWAkyJEKFZVnL
1duVnIHOQYquZnHtoNYSHM3WCk7XcY9n5U8NWbVBhgZl566QmZAOVf4eTG6Gt0aeIftz/kNYMVr+
qD7vlVFUe8BzwxQBJcwVtAHtChhYYyMokXJRtMWkuwsoRTqVRgCbUN+uNO+pStfY0IvdCFugoQaY
DUJUI5ycci7eZjQ3toIvfudkHnNduekoPXXooDTTkqGotSTd5JneT+V6aLmHk/P3LlZyA2PqEq9b
H8WYPSv1ZOU6/cgHlT1+nC8QIFz1oj05doaxDrejjCR7eYync0rBlNpfsvlBr6blSfdrp9TUPIYV
lq0DurPtTV7IobrPkC+AlT11jSoA+5HWFHmcg0YsAbcqwgtQN4wIH3uKlp9G8mDVKySRLv9BxUnc
EKjRiyxTERJ2kka+t6T3Ivc6vysQtvkWuHakEtJxpBtdVWxEGLWMY07wqHYgOp9pm06bKw+k8ISC
x4SmUbq5hYyM87Rs3VbT0H9so6eh4gu0jQAEgmqWXfXb+MSEh4TPRZ0RuFEUYmcTd3xFwN7JOnC1
ZK3KMLoBm9xo9jwn4Z3vZZf/DvtXZGJlq/232oFXZD5c1r3NWvKe1+jsQn10BDT6+mjx5MTx9rp6
hMhDdeFNGlDN1mE6C82qYnCvfcQB5TZ+y0rPFG9aHayXV4XZQrj4JEMcvT1EmxOb+UWMIAiNtqc3
ad+uDf57LvCIgC56Qm65ugUoPkfC0cDmjuaojPyBPd6NcJCEH3syojQWzm26EEQPpW0Lq/I6RA8g
IwhsAkn0tZknMGRqJPkhwbhs2hPcc2gHAHDwjoYaEiDOGiZ8C4W1WhpI46tf/2Ju8FrU4XJ//rzu
lKjqUyvTGb/RNF+IrURJkxcylqqZKTbbiDzu2lypelIct0H1eK9hwPCQxIo/4bH7WrCPb0BJ43iH
euCpGONqDL3dFo+XhyZRukrY0WVi9Zc9zurROELTKkYy2MPyrkwaoUaZd0Nd7W1kzmAsHKVr0Oyo
6umXqqFwBDcDtPn/YEs139t/xlKmmTMF0z+s9Qh0am5L5YJv97tby5s1G6ShH1tThD2TV54Ql2PG
Em0qE9kzrXmkgDfoX4t5CIjC6GNznsUc3nM75qzgNhRMeGAtQDvxhTktyUtevzS7MhGU8h9xlOeO
4We1h+xt/DHzvbtjTzeLKAJLZ5pljCtoG0tvqJq5sflR1qC9H9+hlhMiaHLsfQTSvL+211Zpz0kU
JREzwDWNG00eQCtjXqkvBDOOgGneI+x76DDHzX0ynC1OUDhf9vsZv4nHM4sBoC7Dqqnysc7/0piM
i9FhecVG7OcSO1gkz6QHanjgQWaQmJz98RJFmsY8XQi1mlB70eQH9pEdW8ZT0/QtJ4DCg2sasaj0
xXddLs95x9Onu0wOUXfLFlldhSfPW2vau2m7Au/q2zAJnLpNvr/F1Y1d60bqF2NWZ3iKkI+Z3csG
9yahfmhf4HVPK6HpWW5ydf3OnMqKWuJB87+K2+dqhKuAqMoDUgoVKOqNZLA51EEqqgBXlnVKQjnn
hU8tajBfj5JPT4BrDxviwuIIfOCkly1JEAqOJ+Go3iwiHJ3pmfUpW/pLw1JuviAiYhk3QKJcgzvm
zcD/zF3KkcdTim2L32+Ov8H/PPooo/LGS3YoWT7TuhZTo/N+IObdnQN/5uIj1Rom2LtecHIeHAyB
0BJklotXL8qfiZMpaherTHguQQdxXY+5KoTL2mD4aqEJLSdnOlMD6fozXMBF3ypZZQv493+NhxKT
G6YjxUy3roZEdBscS55BuNZZ30ib81WjSrXZ9xhAVGCreE+KmaEYASmklJBjkHTXh6pOrndyimr7
Hqfe5qHNiyg3y2bHX9y7pJwWyFow5K7B/bAtRnG9MZmGk+gzPcOaRoitZq6TO4x48LclbxdC4szw
aUY6lr93BmQB6uYEQ8EbwM2zEiZuqz1kavawEjdUnjoikqs4qXDTccraR1o7fd2q+maXOyrPmbpv
gABX/wl0/BUbd5F9qBhbesSPJ5LT5rj7sbATA0m7cEIWcyacYofz392C79iNGqUekGf68fctrbGv
lcwr4wgbNn69DGeKTOdcPHmykm0KM3kDOTvOEYC72dUcCUJBUrXDdnYgyAhnpoOsvWVXhNTKxZC1
LMm+j3rtX5jbhw6VVga8Hu/L93wZKb17yFbD732f9RuPcROZfYVZgFxFDVgbUdVhgO9ASVQFl1NX
3QpUuZLrU+vcerW8aq4dnQIUhD59rEdfj5hB1r9lXxDTgeYPQJ/wGZkbaChFTwcpAuV5l9n7bmcs
yTtLx04eb7+LSqvTee1c3/wdwQh3xy1TLAkyHs7aUC/zTdiqwSpq1jq+V2qLAdNh5ZYmub2TxpKu
K3V/bs84TytTWC4NB0Kl0uxG9NeUiy8KDqt2V2xse2eQ2V2k1u/h+ou4r8JlFD8AIg8kFH/T/pHs
ICZUGT1pdHelDM9SQ802k1niTIakanEyeFtRc3RDU3jgM5zm+Kco0UQrWm5PJOdOatOikbSxCEQ9
2BPZlVVyY6Nx7uilg7r6ELQMs8JVORCtRdl6oM5Wzo/gLKV0yguk9omp9ZLK/tFQ2N64KINbzHA/
Fx2IgtERxlTr93SBu32dQdxFhYjKO5lJ3Wx2AqX3UDQu989QpGEjWUsBJ5goVv+kByT6AHVfHkJm
wEtP7ooJdmSlophj00qv4tmvNihxQHYLTxvTO/8EViSb6L8L6/ekF/y/PqpXt1jvsTagkqD6kvHP
zPX7gsXBC7JHxfc0pe5BbKKR0lrCoqkjbZUebVyajAh68mSzAnAWajAjDbKuV/AmGkhAJ1svcNMA
BwCD70N7DEOZumUYUVIL2oGWMl8anBvVXnZXHKdhnYaYCBVDcIGI38Ln5Ool709uUz0KQNE+q1AE
SiBvRAIDDquJmMWJXnNEDBHYTvNWwat/KkRSZG0KkmleZJu6jzA0EGv26KXZYScffb/p5wJ3oU0l
fjWaP3BYkDkGggZjuOfe5kKmE+n3jb7V5Y1IKY0ZckKmq8Y2Eo2WTuYSrkiaUn+Shfl/6cP70m7F
xGIdGYBR3GX9dw8I/xKb2ngtUqzIxPAL4xjjRC0ZZSScl7P1RPpJi+8atm+HaiAwy0hIJnARESaO
6v6M0fNWJtMGIU4Mch1iNMwYJxv8fTLqXzHS1hna4KMf6jDikUmfb5yW7w2Z3y7VHO10FAJ8LCJ5
4tTjUlk3+uG0bwrxdnDkGCmJ230pfhNQCWP8Dtgh8cl819h3JkWpSIEjIdRX31tEo4W3Tk8VHOgD
zTAGInCu30+9ntZQh7ngAJ5LLFxlXqgWRIqkiWQRXCUsxXstVAtQgUzG6Ds7fdpLe4JT85AjJwzL
xCOLblwsjlFcrRY4Cx3nrbRg+/zUy/Ff1HJA9O+topuc72qOeIrv7xRm1iRman/E2HSYJto9OSSf
h+eQ2qYwOjJzHIP/0hnoGm7YbmUC4Gj/5aCEaxujWovhibMLMJ362OnMlNdIZlQtcfolXFzqaGxl
mtycWLXUpMT8eprvdtpeDRN2Gd5U3xPsLHRpuCiH3ML6RJUiIchecdyrQ1t7jtNfmaxGDmKclI8J
IQjYG9+jXmseOj34l1MsrAjFuhi+apV0R/mgpjE0SHgl534Bfr8R9l85XjTtJLt07ZjpwxiBDHoT
MEAEbl3R+6xEqb0EYpZ63VmsxXBtiDOxV20+pDO5eGHCBG90WL3zf343NSH7F//AqdSd8SH/9uYh
hsTG/eR3xQhpSTBnYRy+WvgbfafSxNlmigjTm/7uHtIpR6KZns0FGfWicElIi4VGlERzxb/PE/74
hggxzA0ZSG0S4mguL0pcJUFjLmRx4gmfA3PQyDRHcGGvjBq3r/yxzJUeG4IIlL23YuroBV2I+t1r
E8jT5FK/mI+wYw5kHLeGRwxXWSpB/431XBNi/sUfRnfMkch7q687RG6C8ov96LypyZjtDGm+k6rs
ppBNMWwww1YIk50ZtvRvoD4BKDAnyPC5TQxxvzEjg6yBZhomb7fMpw4zPJslFONRmAOAuTSLNCIW
cT07jvz5PZquwxFjMPiiT92KFnoJfq3zOhElZFzNC3/ECXA4lLII8EdhqhwGZEerwFXotpT2Bkz5
jmefCw5cTNNZfmBvJtcrkEP8thxyQjk8fZYWZmmT/EtQccOnJi0Vnvm/g06syUxMsKr0nEnfGhVC
gVOvBf80sdFkGOvY7quWr8/Em3Wlkazl2FsvUx7v29wza1ndoFOo+S+Msuzd1MjOLS2fTqddOn63
pT9l4nV+Ykhq1ZX1JgGObIDlpoPVn7t1H6pua0HjqPjoptTOCW/zrYhLuP6KUZR5tpuuboyljgwZ
jJ7/ZPXgrS4Q/1j8lZ83zC5q2ZUuTsCD0CLV/PR9IIgLFtfdkNyYt92X4hzVpjZ5eQ2Ct4XG03Bw
/xtKpu+QQwe+UDyxnhQIxTd9K9mRfC/OpcuPGf8OQ6OIafAOYU/gjqhS1TpOiyyYls0b13Y04hA6
jP9orF0ZiaW60EwYBvnY/8mATCD+pp6CPgshRGSOVdY23urY+otfXqxYCevK4xwakEuIllvR4w+Q
k5UyuBD+uW/vfJTEyvkUMXODgtIC9Z/HUm8lFlrVxpcVkFKGb3Pid6HY3auyjXuuV9PC23TmmBvk
Rq6jhIwLye/UAW7U6bkRJEj+YGb5HR5rCHKnXiqAguf12+yCCm1biMJsO9n1ldKOO3E0ZDYyxF6p
4y3zdvBPCo64ms/0WsCkqCKvBlvEM1XPT2bzRbwRJQoWZF3Vod/LAI5EidXy+a47gf/O1Q4w2UH6
fmdZPkpZD1LWFIIWz7+VijWiev/sNRSujoBg7RYUkSPh6KXG9r3iaTSdmYqyZXxBesFmRzIjpa7P
Z780vUC7yUOgkNvhjbE5un22ZqvnSAgSZwY+os8dXX8ghH2WjHN69Z8FwJv3NsLek3kRFAk6g5xD
aJjMaQfiD0e8tTqs7mKrSfrxZ4Wa6wzccT5/fBwG4L9U+OqwIQ20axz2PbAHpp9SUqiuIYTYQNiW
Y4Oq46ofPJ9KvmQLcPAIFr87dgkIES+brXOCOTRI7WW76OgutAObUvUU4QjI5XNyNwSaP4Wi3ANI
CEScAAbv9V9/lgKLLxZR5TxUhVbOLW4TIoGAq6VuA93C8TQb/1ZhPK4fpA1XVHFDON1srDTXOFFY
3loQ7qMJ5qegygTXd8vQRPXMF4dTH0zuIdqOH/g7RgPpSqAqFf3ZB7GQe5ViwSOPGTAF7HfZz086
OeNbjfJA9G3QxF3oNg969nSUI8RY9WTc1WRfhSgZkkfQiOCulQTiVcyZHhuLPGUWpv76sfZJhK52
ZBD4yGKYhAB0FpyRWvde8klExR7+sHG76hj1w83+BT7jG83M8q73iP4wfke/3JePXeZlc4/eaEsG
bfJSeXV2PTbIdV0m1HvDwYdNnPjfjZ2GbMv7vW+otlViDChBuPTDT9cpoqxdYkhCtfbpAPB13eqZ
MKhGRIiD2mNpsvwuDSt4WnTk6DufZU5c+4aXGpVfNzxGReALU2XaC/G5v+N0arje7p5WvMyXo8Gc
rlbuIwB77xamwZmzbrrJ+T3WUnk1RElCZ5agHNLfrrhiK9k4w9Zvxos2eQTuNVRD1kbfd28D4KHb
NmZrV7ZlkXB0kiPLzrughdrR1v6ObKyS7u7/93iKwikaJfBy5jEhak6hFdEbtgodX2Rzi1ILVXIG
iryk/cSgXg8yhnu5lF7HxbBWzwft0Jz0vnhAg0iYH6v7E4GA9L99n3HQfuqZwXJ+T+km9hOG7ddi
ngqICYBxewfvGCWj0+8YhakcjDFlh1vQCnR5ndSgkHsxXB4jzEeKrf32uLGcaq+ifznkqSdCLO+7
8Y8wLMMDVQNPzrAIKsy6YMK52c7lR7TLYp4atWuJvSV7W7G71WU09K2kSZaIUKxffu/Ogw6Hilcy
VVkYUoRNvV7hXsW9DHzxuSifevfpvQIBrA000EMRWD+DKG+jdMI9YSKpoNrSjX7uCvnfx6yDopKV
wVeLdNHM7glnNnZdI+Ie1xmaQVGS+47BKLQ+HszJYNHTN2tYozm//eAH5zhpPqJGW/MVt75WyDqe
iYwFQ3khkQHU3y4OL5h4GxUn3XWp+GxgQmSdM/F44eTyb5xRQtdlxOuyhvK6JcY8hMpxzpn9/PeH
ymgZmpaDp0KltYOjc3Ti0eQxh7veVsLZtSwGUCnM92vBBCfs0Aa5jXDiyKfnnmXC3KTBZU/VHM5w
JKQ9nKJqhdKnicrI14NnU4ASsh2qcZJKLxE+z5eDmbDhqpdXDfXQNBZKpmXWHFHjiZh8OzoFhRp2
3AO/CGGPQv5AnOhpwGm/SlncdiXhgFe3KMvbS0sepxRi72aBQfEjqLnpioi61bEUCX7fQcHroD79
XxQ0Msnbn4KYMhC0wHkLQ2WG3YmbHMaBSkvArgHqJEvgUuduqr1KUuupsfYOChUdjye74ae1HRTS
UlvWYyp0nBSMIBGYmssinkmLb2vi2fKm1zdh5WbjU/XQub9Uym0tD5Eko8zJtWa6ANaJKz59kV+B
AmDWIUR2apTXdhPmZQDykcJq9K4WuzqyWf1uhqD/7YmGY3l8j+j+WuTmiZ7fzUJSm6JaGgxsl6PA
n3Ut/xZ6fci8EbJzP9FOrtWXNZ/WEGoOUWLxC2VsxCMkDPriE0AYiKCWzJqyg7KmfAdnV3882Ud+
pmk9utyonGrvh9DVC8sQakAtgE0PhqtZaGf5f/dXoQbFsnJzBTjKYAiK00w9R0dJ2gZMDnBh2EFz
j8TFzOeQtXtC4qPfOO7vwqBC18axQbE0DbOUO7DG8BfE85eA4gNzzGUlda+KVvWbwxsqKT4iRPK2
SVKQgOKBSt2vSsCPaYA3W4EatvZjP/BQ5Mkm4BF2PgLfBT44d5WxKgUtFWCaAwjhtHu19Tlf+Evf
c/On9n2sinVsXK7rXQhuW6fiKAF4/uKThSlTEsshFsS0U7V/zxzw0YdTJales1kCfKEmuB42dH5y
VFRtEhIn1z6n+xpBuZjJaGkqsoqEFMj/P1sOsVLuMTxo4S7FyidwO15h7PZC4NsqM3YknN8TeKp6
liBW86+cSgWSr/ZQ2jFIi9m9Y0PD/IH4jEc8FC8nm8Zv73UsLwuNbv63XE4EI372dp+MU43EV074
Wb1UaQVBV3dgoryEeX6BoRd9VjmTVsrPUutPqcxI4Vkiuo2UUtE/FurYDT2OOExAZw2OeWhLE9dS
FBVgmxvZckAbr7A+hz3iG4dgP0/wC45v3hnsaoY3orvTWGV6Fy5A90vuLddC7DSpUuIYuRVwtln6
U+xe6u8ueIZiXuTGl8h3JuRZdM1K44qGHZxrLl/Do7zo9rvjDe+PksTyWwje6pevniyGuDn1rcb1
EiGfu2IbICuUGCe0QzWLXvovKiwyBqrtQsxiQAqOacmOAkeR9ojIjsa3GnrFfFisQekof/V1llhw
UbotgC8hWLg5/+RHqwXMfHa7ZIsiLf7pR8sBNn+h2x7lgODQsIALjmOuSCclC/rQYh+MRWY0Ncwm
FdxaQEVS7TY2bNg0gmBAgeHXC9y8GFkCzdwltVelaqsEx/ITbF+f3fEbxiZ+HZVESJvdiNEDGaAY
IWGhm0Y9AE3G0O+CmqQfgzyGNBCYueRFdN3OD/E/Dg9Qizyb077kSHwlgbCaet4A79uel7WH7xlu
SjXB/vu19OApoa0f8ItS3knxH4CoGACbKb/+I3TEQLDxT3bCdPce6EXwE/JbK/x47+6VC61ndkQS
osILvrm5+4xjLwahzlxL41n5TL4/i4ow125pDhsHcbfKqZq4tEPlYT8Q3wHxxFmwKLTxG+o6sADU
cFaIjfW2CVclOxul/G3+aADK/Rn0T8Ij2DpqLknkyAJ1KppRjO2jV4nsjKXWo1QZ+NqYDg+2smQ8
H7RGuAUo2ZgOKoi0lKf2bjA0xQp5Ho/VaphBpyIcf7EjiEQSajrI/72Vup+cjDUeN23yoz0u/47a
BYw7W5MvlX+VJcIEm0dPuJ4yyGpdmzIm4AEW0lLdNQ/o/9WxK9eQI1T0Fu/907FikPx1uZ8vGu2A
xPuyPnaJSKv/3iS+bPoUy1rxYP/70oYwQk92iJQgzqzgPprDvE9VYgs6EndlPOt/mEFuCAqE1oLw
0Ai0LCp3sTGgfCWmwSUZLPjKvTz3w9majTl6iu1BcYaVkb7InUgrPoq1c83Q0XGWbpTm3fD9BSdF
t+d1vK3foi3zDOaBuiNjiHQNk2Oj9qN0AnR/Sk6TXmn3VXvPytATH+HLYEEJNIdsjH3SRAkRf0di
MpuGu0rP9eMLixif1vunHTwYjoEcVudglONDWyI1OyGqEAcjYhLL/ZbjT9Ltd23wUSMLoELY12Uc
aJqgcpwKQoECdsGTdUc7WlO2dnGdhQxKVsGcK+l28rpx31WjdIJc7TEOsXIbXWi0Qw/7aBzDNuwA
rBkrAmnaF7NFSu4xaDSAVnJWQL/6EIn858GA+R4qP1nN5NNJB2VlB6n8PiD4iCuxqL/1Cl+FqCBX
SvRaeUX5T7dCdRLXUf/989uYLmGcPpmEWFcBsl5PipnC7VCKHyuHKumwaoMh2DJN4V/YOhS2FUB9
PEEs7UtrukhbC9Sc11k4DdQFhluTdsmA5D+Pi8e7NKoeMHXVocVKRUReHGpgV+h0WpNXACM6Jlji
zUUAqQ5Q1z3q+WiXJdccXNxmU7nF2Z/X2D5yzv9I3e/i+LzDwDx2eFvJZCthvB1D3rdAkSqU6JnA
KD5W8BLiHxyW+V2FasE/neR+RPZ9BcX5jwO7Ci0i8XYoUjjKoI21T/pRYSVYpU6/jIW7FoWVwwh5
rCwBuqLYZ/p5GW2LH9EP6WoMf+dRoyvxYVJznTCQh2fsWQdB5Mgu1twGNkur0NNAk7E/0HdTasT7
Icd7gXcksse4qut5SYuLygOzCXK0+6Q15gFxZodVq/C1VeGABmYpvD9ton3xJDybglfj6ghhFBrd
AQoUCF27Swl882yAY8cK+6F3XGQu2oarGw7zUwlkKA/D/LroFcUm6A+5He7rYp7Vgi9k32iGsrwT
gaZUh/5gzCDL75I1ypPfPAly6OlQ8OaFUNzgSSzyLCri16w3VXIj3sBaICY8FO9bpjH7j66bPZzi
DUMvhvs7R66rFIlCcKdBGnGtGwcpYMBIOCp86rHNtOsrHqPaS1g2gGgHZcSnj5Ca+CC9w5pRmKjA
u9jgKwBHHxevEwym6mHJ/MTqh/SUo2aRbr/wg9j20WJvm1XWCAH6g9tmkyr3OGht0TqL5yDt5ZB/
rqtP9qgNK486QN8nVVqzOUw8mPpe7G6LskB64898q/Lk/zGr9snoAZl/JLa2ClAdjlluimqGAUZ5
Z0jWuJnJmSHVlFQn/sUx2OwrmgertyLxrxdeFF8wiqJu4gZNzRt6FzIew2zfton1NOr1jLDjvDjB
6dZKClMnyipvubXd+uagyEcMuj9LT5SCSV4REePPiM2ugfs1eBFHhQExKLrgtHZyB6p8T0/o4G3F
ibbjoxNhbOq/JuTGvXr73FnsCDCAnKlmf5Zfk4MttQO5pk7Ax88lLCH+bVB0SWznDeaIlUyKOhnk
wPOO0FXELI6LDFQ42seifkiNtKzK1G2i4+CQSWAeRZFsWnBfKJxXFCC6PD0DAvMkN7iWOV3ba/hn
AB/InGX0hfBKufps1hXLmFo9iugDequRFnp8z7aC251xf8KT/D00w55I8d5NfymltLnMHDwy8Rbq
oHXJfazuotQ08ezSZI5+n20b3Awu1MyTy/SX9x7Vwwf7SwHrY8WfPLmEpwDefKXWf2bF6kGpuvFj
4OdeiwcuO0PaqMUBHGWd6WrQag7FX49ZRytL6vPdUl5Hzko59AIcItIwILVnvEU5TUjmDVCti0XC
wEJZFuVoUGExQ6IWYQcN0EaYMrsOXeOlZ++sUXfF3vefBmEdLfrEHs9BbHkck5sPbd0bH1RBwL8w
AnIvRk7eN2xYmPm4Wjp3ET1sq/lYHZpSqZc+kSO78dkjrHKJmlCBdcMioWMDkDr1HtU2te27SWBT
u/gOP/fiBRAU80+QMtVRRGN+3bkDQAAw1DnYxVqLjTuhnx/l2GI+BpSOqpQdzx3mRifVOWL2T8XJ
b39LBW9KR+bPVhLxY1nPeIm5TBhiupG88zx/4PZSA8hq0cYcm7uS0DHLcXoP9rrdJgF5ZqyGluYq
rY+uDaw+wQ8/kEna6Zw16plm8DaaL/YkY7V0wF7SeTeOWssOM5PMyOK5K7tcwHnp+1hgzJ++aP/2
u1BCXGSXNLpoKbYTHYSr9/E5NTfWlbtyKVgZooUFZO1C/2WwQsMRQVT5p8eSp20F1Bz3WxsiruDz
UbO36WQJitfDos2DH7HPo+acUhcvRWR6abYp5QiH+3P2+h7gOKznTVAB/RXVpTdii59Pax/25sAV
EHh4tA2dCE/LyZlenmwYBhzrmqefy9pvTEeiU04zPHlDFPUuYAVl5GsNG+bpEnUPC54/585iA2eE
XTZ3AA2KhofaJ3AbPbqkb4KcNeNxYPDp6xRfmAjTEEOKMenTqfQbXBCBqrHbKvt2V4UH8dzbp7+/
kpL3ZDsAEnPUHN0IKD5ZJSab2dZIvWBhlbSV9PdNwFwRqb367zKi8V+95T678pREnIXRhU66etuS
D596bttzOJTATh0hmK2xvShx9+tmww3PBns67xxNTkN4tt9pHLsAPeKALlQMubz2nJdvQaYdHOdm
iPuxARgVfoz+x2gx4iH1d6VFhvq1YBVGMpPgZZ5Ob36cVNB5AvZ/Xsj+WaTJLiO40ow5iTy9ABop
YbAN5UKphq98kIh6Y6WH9Z8ihLvtmvlQTDlQ+2Lql8YN3IOFtdYYZ4Z7vlPkhepJzkfRa0WfTifq
iEugSAa1glZGG1AVBptEcg4taXhxXeekOjOPJ63l6bA4vJT7Ab7diDBS1ld1IyJOm/arF0BxqjBE
DiKBvCyAsDqu4mdZHYkb9elIQg4I4HI06XfKqsVDAE0D7iY8h/Zs1hjbjKB4IEpKlt9XRGcWZzD0
2qoiLMfF66bfALufSziM6dW9udwejcvS2j1Fb/g2hg0cAduk0mmw4k1AtrO/GlhWjv+PgceS1+KR
/zx40b66lEBXYQblkLb/8ylO2IbDHBlEjuvYrEiAz4y8TGnZ8ptrj6lTE7ILq9wMklgE8WzeG12s
etz7rRdcJVOq47Bt/Rh6fi0WuumLMEEc8S3fYoJWJRpYPCqFy6Fi5XIt1IXAIvjuUefRcbKFAP4i
srcveAJK1o4/87R/iVwbEDnTZPnlWtFXILasG4oIIAshQupzupm7KkixCmv6SHknvIR/lA37bJn7
ERy7iSbyFhmw8WO5FbWPvUB84rLeu6mkN1LZBrWTga04gGAwdkhX9m41xTC1D37MDjKQTK4pvx9g
tyaegcvvFejYz+ZvK393vdQbH8c8MP0p4PfD7ldBKeWzNQWK05eiZUN9x+n3Hjc9B9fAyevMLAIE
ls1M+Ep0RZ66wWFsAb2w6avZobEiqVnKcY85aY66bWSVkyDSuT/Od1ZV7Yh0BwyBq7Mbwl0NtCSj
hFdzP9Xq8LkLCAjMJeZmnaLEew291Ye4ZYIsk3UgEDN5YFn+Uz00lJwRUWTtqN2/QjbElIOAvnQF
iDn/6Mba8WliRIqDiL0Kn8Pu2ALl6Q2IRJ3M7nZCC7fOeXjAyGNZBOaHNbmtVmZvLiMtJ2wtgQlH
2e/5rjHesOFCm9leFk9JMOV40+m4RtxCYTd59QQLGN2raqw6uyu2q5GHlyGHkczSvmjzEfIhr4R4
DUiWtYCTrt7gvlXigPQHmtJBsMDTGDGjUjMD3AJvNMBMdMIZ2P3VTnJZerqkwcHkLuBZ/U2Psb53
dgjPke4YxISDeaRUgyN4sZKa6JRQpxqol8hVlfuKPo5HoiudlStH11/G1UF+vUzYDFKPh5tzTBjB
MGfQElY8nDDBIRsZgYPHyOexn26f3JfW8CSm2M59awFb6gktyG+fwx9NtW9GNlddJ4tubowl8dhj
IT16M8FPwjyYtYzSal4LsCG1iq8WKFDmUpt/o06iEAeEoUDOcMWV45mKSt9ZzUsgCxSoZTCxCY+w
QneyKTsEFP/rRdJ7a3xRcuStKDuiI/QvzTV0fO8vEmmUYq7/mzPeRwjp0xUMBQnJwFCPPDmFPnBZ
0Mzo6/Rq08qiNSOFZzasBybbtdbSAk9WuCvBHlMbAfYilHNbUIkNMqPn/qCOpgBYRTh/TgWwHB19
l61XScJ/KoNRUEo4MSvJ35AXB1lHq4tchQ8eg6rxJv+VNWMi6EOSBT10cWpvH+WgxfYBHOvRo+Az
DYW/mUOuWLZbtvzdyLCwHp4tFLVhWc2ZyWuCA5/F6qzk6vmwcx7DLm5qPf1u+zfaPkKUJRoKGW+y
6xGzazzCwTWGZBvXfuNfqwwXZZ2xd64BNtFXzuV1Mz0gq7zDkAfw7DxG0N5ucWy0scsoXvEltWEm
xVX6fw87SB3w9MMJ0ONUvUnhfp7YZyC8gIgwM/WccEZVC5mbN/L4sv/nhdkUUR4+iMFCsLGNPbjN
fQMDKZAcAqPKQuklbKAq81PFmNuoLIlh7pMbbLcmT4pY62KRour70A5+/MFXhGRXkxh8vT48W0yQ
wG16NbYQBAtXGb6rUY9qaqn1AN34Y8Y95EN3p56yf8yZwGf0vQx73jckoW11HJ0MgUsQRMTfzvxJ
6IODahdq79hMGSezAmIqolo2p+8DZ+Y23msxNR88sL/XBxBxdEJHRKsb2tt5CydGf/EXCSGXQJqq
BCw3TeXQQrGg6QAwyIIc1wYktlaRPjx0cUMMSqdn0NPuzTf/g2OLbCffjpQogzdprvueXrjDk8jK
sRJ1bCV9s672+09rZSlUv0TNlyYPyEdRPnuPY4Sa8oJNbhuaSoTl2vl7plgKejqNweQas5jVvDlc
9dsv0qK9CHyDVResLapQOKWIJeLdk9pLkpAteKTE0zlGB29JFbhfCpKQX+Ju6Eo0/kVEGWmT6AW2
ge/lYpjmhG4cPMSH3sQQcfoiCKF63bA1Jlo23zfbDYyfKl77qhLU40PqQLzKOpzkNZe54cnZdoqV
ItMup0MTmOram7y98GRpN3w6xT9OCe00g2Zgb7OEj5qlZgrTlLFh+1PKMhx78djInaF8j0a3RTd8
J6CW60RD2857Mh2qOzJV+mHpbVLgNueBVKTgkLDov4nQbtM+FQ/ijYIi+MQRXBavdr67EYJ5EWgu
1yY3NjooiCGTfJxM1NEZOWkphk+Lj8kHlPo/56fjUiCuSO8x23InN55Q59YzUl+XdWd78VEEVsKT
5CIKLbkmXnogxTx8g0yS5f1lfDT6qtiwaIfUSuzComEXmobawFC99jhW640POHGwT7IbJaA1Ts0d
tFdDy69c+HLJ8gQqaNEfaIRQtm7BSuARRiOmU+JgbVI7RjCXgAoKHgJG2LcjOQsmLLJDQEKaM37M
rw9V7fbx4mFFBth66CZV0QbJfHJE0ixW8T53u/XQaTA2nC7g325WU8y5Uea2JMY3olXkOXtaMfCX
e5ZSVXukFr2DfxUBsNsl2avh3q+QjZP3cUrjaDGumR/MW/QQinPzyRe2p1/+AaU9JjVQs3FH2cip
iXBSFHqUzQN5eMVql5jv6Z1EQxT/I8OmX+a7Dit2S5LhEELC5cGonf7KJz62iv8nccWJQ59j100A
qvlB2g8ru54EMXKjiF1oGIU1N1WGZhdNuaVGmmXZKhd2pAEGaMRtOKciAWfF7tTvn+DDEEfKfWES
MF86bURqiZ0z0IkMxAH7BMVrEWGiKFAtXigMrxeoboRebR2UKWFyXbRVxil+TJLBqNEQjDqCHnOq
HaX3FvDK6+wDtuRrgpRgqPjR0VJIFpyfAHz1Nv7G+P+JDMwdlGTK9+Wlxlx0ROYlhmcgBYUb0b+X
Di1PVv+Sz3we4izFAbpMYJ+eha8pKohl7rkR5YJFY7l2P85LSq+1H9zGSQMbNZxTSAogBxFGiS3o
i2HeJMf996rKG83fFG64s6iDjYCOCeR2Jncc0v6+/dCAEba96+eaAY5ZUXuEX3XBeabyRXgLPN2F
qj1P0f6sBKkRqztCSlhHkH6pRJjdXbFmffpWWb1kVPR/QW0IbnGnUZbmX+9NX6XT7SU1xc7380fr
4MJK7pc94e/4NZmftKMh7EtNjW+i2sqtIxc7Ui2CVpBUNhcRgoLVI6/ghm5/vh1J7WZ2ahThVO5e
11Bz9AbbnL9UyNAE+Yu3vflTH4evhXbMnPKuN97anBGbLYbI4nTHwPoLu7Y7wJ9Ve+A634sHgCQs
J8t6dipXYfUF8yMcsISicIqSW/NA4u6TLQiOxwDIZETQcV4LqAIUAbdcpTgK6J7lJ579kft0+9IJ
DX4YnvAza0DycRYVKyd29a1ISzfoAVF7UT6GiggrXliHo370wZ3cA9W3PfhOq2LSAQxyRxfg69Q4
mc2rqZ7CFtkw2+zkrT9Mo0O05tq6qPoUb57MqC/oJ7NhvJxlfCMLX5o/3ic28ZEHRsdvMEqNEb8I
vqW85l8cZtUj7F6MLogEUGMq3LaO4hvuhW7hV/IIBDvdvg9/HpqOmOTKUIkqLZR4Yv1vOH12GYKR
OH7LJbI7oj5gKbeQVITSMkc/Yi6SOGdnCd/upo5sjltSmnI5irqGeiShqxZPzIaAQgqTtRU4t+07
2dfwg079mh2yM/K6BZYmKZasjnak6rXo5vmO0FPnXl1jwRjGUw5/MOvOUXzbSB/8g7K5kGmwGrba
Xo7qPliEzTQgHGyqpA1xi5Dak1p7LOjVqtd0cGIqVqZ9mmWxHUWGYf+ebhe/5Xy4iVDS5J1lfmsN
gZXRVYXyJqhzUcxJW3q5fdUZ3Ocn4krBZJoU1qMogB5d0omzd/omkw9BSi5/stVKvI93FMaQvPZw
6QhPdQqYPftbLYqKjlkflihg92QvlFKN85OByhRlllZ1MWBTO/D1hEFLO1DmTFH0x9QB3vwAWh9i
P7zysIQzezMe5AArvouRfm8HIwHLIcWcjts+gR9ugLoqVQlHmcWcHAOplVsEUcW9l+YfQvsrzoei
vkl2rIaOVEzXWcNei7DPRxZrOnFt/+jVCNXHiTeSO0nyhCTHTzh4lj3zOJftUB23OliGsoqxZM8i
74byPTJFXz4X4lKsBpmULd/kcwbHCFZuU/Xsyf+Kr2jWnKst+m9XuXJJjlEPImUWy5nVXubCiAaW
b5ElLeW7kpDtJK1qrF8B68L0a8vpPq/0wqUMghZNb2I+h3/8hHvWCS46QtSgyezd9j6mrnD4K5JW
oxwLZBi+3ikt18Hx6bBnkxmWd6MwVeW+D8xcZZ/Odqj67lm/fU858XzOMNjmI1H4Acx2PBuf3NLh
s698bSYazllz53Xi1f1kyuElHtbTvmteGImp88CX+0qlymBixPNjoDWgSYrc6Sx2/WgEgXq6PorR
VepI9d4tyzdS1PvoVCyAKHwIrGFUQnCheaq7Eyxnzsy8MBTGEJzNbb1eAa4MNuQbpyetBzPum0a4
PUm9kdM5yOG9DdQ+HX0AroCZSTAwL1PMF2F10z+HwTeslnlcuJHHTgeHr634dybUYvlyDNpJlt98
oWp08ZmJ32TE07GG/2WzTqznZAFkY+2hw4sNpo4KFBN0Ko8rAxGQoGYH1va+QJ50AWuy2RZLeluc
0CAr2Zjvve9BcvvX88cSuxDjxNjWTmuNun7DTNBEGDgY4JlqKzCtDRAKKILzyLvszrqtSPDePZWs
J3Nva1VAXCuVEK7FB0DpFan2QEsYlR9QsCUYcjlhxpmSBk0U8OUJfW7k4Q7HQwa09N+pdQ/EkNoK
9O3Lvy4ggzx9IJaAenW3P8yPmznkcdktqhb3hFzIczRoAv41nIdma8ogGh4hfdnVLqYiAvbkEhp9
8wNQLPUsK4johztsUNS+Urt4mZcVq8cKbsUod5Fu/IzBz+Duu1PT/hAlfMxncqX1AobKnJOxlmd2
QSeBUE5gRjeve3/eYANq0IbNmLkoxX+fR2ZDp755e/epvRzMV74hsmAXsHjdxDvImHhNEKKRhvZ6
aFmP75RU7DQ8nb7nZmp9vkdtCgX6072br6cV2uxtXMq3umc7YR1rqp+rz8++SDGcwyl73mKOQQ2m
iE015e5AV3U33V1+ZijeaWL828nWH72MH9YvREMwnzlsyiLWm7tX/lESLt58Ys8izmMS5yd5lS6O
WalXFIxBnMGrlP51gUdCf0ftORcN/lBk9SMjRhkSL8WYUiGLLghwlOpnXhpwE8zwPWhkwzEY1YtI
6JiwIvNhp13/LfBHNAy90iAHMvKGmvXXA5hJzUZkk0K+7aUQqK9NdL/zPeH3B0eD4vkSopJLnLKD
opJRbSDqLrfghMmHlTbg5Otm/D95N9GnWxhitZPK6muK0V7OB/j7cIP4vSQICaCfJTSOWAywfpMQ
l/JME5dmxgvmKbX3lMQCBctxxddiyx9XJARX/9oOKn/aqSJz2V+Aqr08EbIYWSPI+lowijELC9Gs
Z1K2+45Ao6MsrCUzuwaeiXDp7w4vFFpY6MhVYcNGv0/XELGIt1aD6nXz4aNMkhf5OGduxR1CRMuT
TZlqVc5jAcr+AL1dU/kZsKd1lgxT4+I4l4gRfjgGoaqVpjlA6mjyuOLAe2zc5or6L33j6yN0Hf62
aIs+69QTAohrvG7NbzyIuOCbsMMK5qJhjTWMX3VAStNPzQn88ZJdX1VsqLjPnMYBg0GgOKUIZdbW
iJ0mI3CUaYE+zRv+Ts8ogAjHXjRW1T43mIJCxJ9eH2JXaG8YHyN8eseayYDpvLsIQz9A4/dNA068
HwZtO84OYuqyf6FiIpTJoaXQOmhXhsim2TlSgBQKIKZ+61LRA7eg1dxEIuCex91xA0izg/JgskpI
24iro1zacOjTprOLvNoDpv05/MmvvasqDsnRfksLAaEb8kcx2BDw1pn0WKkyNkAcg6rzjdR0+MMT
crRy+3xj2l2asAlZp/FicvnZMMfDuP7k9PG/UdCHBwb8D0I1dj7H+a4BDYywVT9TVJIL7n+nVOn1
SZG1xwwxMRirolMDJzPCnrfMp9v8wLJt2bEQVHAlsJbtOawR2FSpKlKnmhwn1qzbFogZ8ykslotB
NY+Ix5jUVbB/7oJEhb5dRmN5sHvYD0zjg9oT1msdQoEp4/x3Vxk8LTJbQVtG7rzWyT6s5cw10SFb
qvo5bXyb63K6dJgHT9jerv4ylNre2L4iGlRpnQ3jTjIueYL7e4QFSmoo2xgm9d6hXhYBDQ407byr
zmQxAiRVSx5YfhEQIXsdmww0nRki97YU0YCy5pGSfY8+5oVvmZt0HEgdbWuk+prKul/Ynm4efg6g
pjtlQ460SSwjbhaTWKXCLGBWyWBfefQUZXT0JuH25cIJi6ScLz1pkc+yn6VAgILvNCCSm13S2oXW
2h8animwEi+DKjs+KgXoPk2c5vP4XM+a2QDmpvwqr2rua6yeFS7GvShZB6Inue1HdKLpy/1/lj3F
4bJejaG33JSYgTYw57nFvfmh6z+2FScwKXghXACmD9MHSOXBZYmNE1gtEDEkhlZ93BRJWrYuN0nw
6CTqsTMDJprqQBdADuUeaXWGqzFtwDXosJrieotKvIticL29TurDkdN2Gt0un6x4QLyw8fSd84Uk
r2gamXasG08x9U4B1RsNWlVU3NWxq7edUkJzpJ1Q4qjRgL1hEzDyH1hR7O1AHIugWJzfMeBZHs+G
rfCM4zXalUUHx4OMtiWcslRve9NnLLcKHYKXbBUOpubxw9Uuu6B5bfYeLd5zlm4ktl+dQAFHUvhk
Ga8N/nlkpnLz5x8FVsM0qF3cxggBmRZN2DJsokCfyDlcEvLTgyy2meyWtxZwi0ggM6uKmKCp9BnU
QV8a8G+AnOSHPV5LCP8yJff+1kFZHi9MVApywHbqYlyIsrKWkTzIlj81muRv3gYGATVDyfl6tSod
mDFcXv3gEusaRmI1qv4SB/nJ/9CnHg6dpfRiQMMOr1JUTaq3mU9w6HO+peCg3C//8WH3GfxRuKPp
QcRngqpcd3jeqIse4qs7fg9iejZmoR8DqqCkKyUNNijTlFrBpJ/8gDgMzFG/9x8fHtanGq9cM1Ve
oChELyPhr4PEnp5A6oayMTXlr8C2T6kJYDm4EXIAGA5NOmuHSAw48dRBrLqzgc/GZEDkzH3lv+Xl
XnIs2LSP93vb0Q7hXLmvENMTVg9LMyOmmOiU+Dn1f5fTEV5aVjuXypg2iK8fFsUCFp6KhuEin537
l05Dmp/9GSYGieUX0I3POg52/Vt8XgvfTK9s3CSMYRoSCDrOLKRvWfv7FbUYMot7yFKpFQUm+Jf1
lcU/y8P4e50tKwnyYvBc/NN6F6ozlXIM8mjgXy4LtYipikAKCSHFdPGBYuPQjG9V8Pme24R8Rxqr
T40bciItp1adTlOAtSc5VMiTbyUuNgvhBnSRqsNS7Fu51Jzy3LRLyyKAntRr60TrsSNCuUHNv/Zs
rIvUZueBbINClDcUgtLt/BU/Bo/XmntXo4EhnLPC6SFCVKeCBNRrTzhY7wT+/QH4cg4cpyKTIkp1
MCsqd6W5Ai7++KXVtXugLTMPMk+CxFFT3mkH9VMRTrh6U2CpCgBjKKIET5iq9fSe1a9TKLIV0WfM
1sZnZokS40J2+qBH3T52W7dllG6dwnrwFt1JXWj8RdmkDI4Y6IKKeJARIwYa5E5ViJsS1jz3Ws0Z
ICYzk8bzN2I75hcqvkCjca/+3gDWeJk+KZXheFMl/iej4ziSe+SioIsB3cQ8uPBkDBlsC0c3U3WK
w+zvlbtF4PVyn7o0IJYKYWllAwNic4B+Dcepf+uY3A6XkBoDjNtxcXNhGNlMcagInHcOSU5Trnuy
Ib5Yjw3H+QBB0H3MbTowq1ug2koOZUFrjgckyYiDp+BpaMWe0LXwAObhYI+XX8g6noRO5VCm2rz1
BuwNZ/YCOfS3SXChf7JEDeT3PQosJhgDgiEywj3BfwL72PuYhoU/qzHakI0XhgSJhoOBxwrJ4QiU
WadE2gDN17UrfOLlO8enSRvL7bQxprMfqZBbiTGXQbsosdeCqw4pRKV7+0Usn8fZXxL/jQTGPAce
gg6HziraHndbwjTtu8bwzPc5WPXnW7rr9w6l+0kqvJ1fEafS8n9Wb554fszYBZeyZKOWBYNcbphx
rzCIEpIGXPYCAu7kfuXNimiiZn/SitrnJ9SImY5juTT67zopgeloMh5OOfglTccKXCAW//43luat
WneajqYBm3YPXjwk9AU9jj3nuzmWOjjDhO6FpixSoD6sndtU7HOUDMOCcIqsMPeHQ/iDgIDFwa64
hY52O2DRBOMXtm6TYrivx3rsQFuCji6p03w28fsgTkzAHjEvAeigGQbxlbRNkENF6IIdNy6IDnR0
io+efZlXp0Re1tjhMs+JzIItTwg9WcJvYMZx357FiW5rDepoNJ9KsW9pZUZFvyBEd9EGtWKMwYZ0
Hj+7du03BwNbBuWDhxw5a6r0Y7sMh+yUG4JiVTQzNjMysEYJwVfASDSoxfpYgePiDmknuPxJ5qXC
0yY14lA6HW3q99A0UpgUmRvim+en4nxp2hQt1LkFbgwLhs+fLNlBdLn+uSkr70CVdLJaw7cKM5sk
55cocjNzekz4INXHT+Sx0c5OzMiGkqqXK19aMg+A4PD4vFV1sMWKNmM/FaF7LtVHoQdmn6AvsTSu
6/JyfJCggwKUo9Dfvu2rxc1gLgn8xAyMuXZCDzI1K85hW4aXdV1iDk9O21UAy4VPHi6y14HlVr1D
pZ2Ek08wsXprGMYEPYiN69I8pJkSpiToScOWjPZ4mXBYlFfXOWRB6E+SuntJYPeD+d9PLcHF6CD8
4hhFpCGO/qJm9IVkvaqdBvs7RSjf2cU8pdvPeAe0/59xqh9qmumMaJl+Ejpw1yKnkvm/7agdq9Hs
l3p2/xO/WI/gNWB5Ox6dgLA6XbSVmAWCxUoRwFf4fLHX8QfoNIWNy+54boByHpThXdbRFcom59h2
9eUoUeWP39Zx6TD/HaIqTJ3GBsbYR/vEUJpTTkQ8QOxV1eVcpqgsDE4Ebtdp+ze/6U9cKAcExaSJ
eb//DovxcCmuiDnbzxLIL5tiaGmkzN0yTvsXNFmcg5yuTqcLnYUqHdUUaebguavxOvxFWdmj9EdY
wq1Blq9yt1Cp2/Z3iaU4jrNnhxAkEkrrEH96dYKFMsOcZZDMdNwMgiHZWyg89wYq4DogqzXfE7Qm
5mB9Zl/0aiQ2mnqaTf93vtot5e2ivy9LXGMbKtKX6Q1lgtLX0NRw9fgojF+6liDZdBR7ZmeyYYNp
eCJlEQ8qZvq6FwJYdALOm9B7ytQVfYwRPS3pKk0A2PfHkRMb825PubHF2usO6DtvpqiePit/NzO2
W83YUzI0IZjIVUk8OfTaSlGAp5eaZeAz4clX6hmciysK1E8iuHw7Es0vLFfif+SrbrgbvmXhej5q
D9ok17ubplEcoQ3xQgCjz/+/YSfg36zAKeK1+dCEQfT27DJQbyitJ6iL/ieMMlC/+Rdj5shMyTgL
K5zo2nrx02FGdE75I1yUrUZ6gnlR5exTD//H4yxDey/1XtLqc5es1ju4GzXKZ5Tck9apll48ueFs
a24lEmPZSoxJPH8RQ7nCMy79igz3kvmmiB5SBl2JwzdSNXxhueSi3b8Di6H+frGESbPiLc4rm14a
ph7hQaWaePt1uAhEr64MVpvcn/iSQNWY+ipqvw3FhyWvwCplE053jcMkmr4sAvhCOXTVGwZArX19
IVyKuQ2GXEnepRNUPgpopEHhJOeo7+I2tTDXrDDu+DrdlrvlEDkJVCyBkTR2w6sRrRPsEV2k3ONM
jkdOmlF7bizlacLQEddYEcugOLi9OXuHBFpU+Kruitl6bxG7V7H8c3EPaxj9otBUGtSvXQQ3if8E
DVKtv0gO3aSLfxdvvqhshTlL5/bECRYxOep3dS4IG/mWPOJuPyJIuW0rS9+8Va4pbPfRkv+n5EQA
miuWlqcFvGBxSNH+3899HUu8K922C218+9p77AhL7ls2BVLAQMRkIaCf9YulB6hBSv3RgsluDOZc
5dQdcaI3uMSa6AdkEzOwjiPZyaJ4DPtx99ElNZLnJp9uapb5kET0E8iy0YLjwuZETo9T3TyJJnNa
Drwwdi7jt9lDedPv70sKhy9MLAEegZRwxjwFVjeR3364fnkkCaAXhGK8pfk5AiD+T3vC+3Jssphq
00ChqRo/0Y+y5UjgxCgtVdmWiUguSnsMm06qtFQqLKpm1rOprofV+QVcgrV9/y2KjuGq2QaAqs7Z
7oJjWUV84auyPxfhJLjRTFCTH7wJw1YucpR34mkUFVIUeDcwe9aG5OomDSasDJY5GSNHr1Yc6+Eg
cm5ichYQlw9812aijFpzXjEVAP5jLm9L7cai7Rpc93er5hF71hFL+gghKjEOlgXB3zM+wzUvfpD4
XKq8Ed0fe5Lpd0YA7acHq4/TVF+lTyAfsTv0WDrdqFnb2j1k8PN2UHI+6Ndm8LLQFjaw8+Z/NP3+
9pRZ+2a6hrQiPVHK5PDkOnCLocXS0uI9moxUZ4U5NpNAKy9dErhAHHEOdG2r4SfAcaLlUmKLSDAA
fiCmWfybfaFtwi35AHuv97Lf0HqJ9zwH94ba9BiaxBIDaCjyFF8Ayns+ysUuxZvN3ifKg8WEiBfA
z5y1q8l1PAH6puuIfF8VBV4ccDS2d1sSJWZv+9lLpOGPMoGuEw9e2DCh3FUFerAbOJ7ilcpo9NhA
BbrUWmsZTRfaV4rYNx2KC0mDhrz8QiNiC+9tJl385cLC1RZLpwrWANbcCkZ6wJdKVEJd6JkQa1k/
6c77udP1IiGOqIQoXY7XH+KRaWgtyHgxGpTk28w/RFPegQ8tVGjaqwLxdjQtGsrMdnWY2UKlAkBI
4AW2JEP+rO/xJTG7bY9x/FH5+LDRpt2wcKUBjHEJWjmP3/iejx3iGChTpfsnf8850N9cvvfjpS1k
mmTxDLh/NUbQPRtqPo4S2TnOTwVrsR2ykccFjrQ1r9eSc4sOW/6Zo7NMYGh95MS+f6EJpvrbZXjU
RuXjR9VNvZEvM7wR/jAdZCS2NcsPGXMArCWh7jWyeWtj3YXt0Y9hZmWxGZbw4jZj9pYJW1jrriY2
9SSjGrEFjgz0bF/t9sWdnaXOWRpVNf5wKJE3rnmr8GMUIPIFRDujGyqQObkZrcdXz877jpH6TJXi
7T6l3JGVOPAUsvffKVaNyuwFo5SoWAYXKjF32WMSl/vKDsLlLEhdtZc0TPgoGZgFkhvj7zvwuEg4
HJbn9GqoAFUiVsLeHiv6g3F6WR+okTFaItmPg1cqMlUi334hkVhT0jsQOXAKCom6vX6WCQUe2AGn
r/MCGOUhzQNMlmuggfBoBICe2wbztrQLQ/r2gVwS9XMTAQEYOtQSOPQ6mtUapGG3xZb8yBPJwYzU
FDyH3z+U/wO3yD2IS7h7+RAdFP2O7TG7qWeLtuZv/WeMy8sYeOWU+wu+1fIv5jOI0gUyzAieWMXQ
xNxRzkJHP1ohwG7eDZWhToZ6vOmwXZ483iylhciG/5MzzsIXKuZv8Wrk9rkyVW2yJ9+KdHWJQI4i
VKNn8VCf7YD/0pcgJtf4Ee6QtiTm0pLuqp3ZORQB4jWZQcNCqvk7UnkpkW0NqcbXbbp3Cfekl0VO
3ILoQZoJl6he1CIkrUD4i4/mRAk470UO8HFoqry9+9C82AtZT//L4X+1OUgBCLvRGg+jNZUhUCgW
jmCfqVr0dOBk7e0LEjMarzBRKomNFkvWraXL8kx6jaXUmpyheYAiDepEXJEXj+yYxHjVlp5tpnVL
FjM6Cc1xUh0vbGcDkyidGP8RCIwAEp7WSCTpVtZ3yPhxAVQLWIge/mNvP7evypaw0M3bfYy1zevM
Lkfwmf5KxLgJls6YfNUorDSknh1/4yqYg/l4RjnyFO23BqgSiyF1UFSGqYwvCoXa8m0jyFgJTfG/
w1Sq97eJ0vVdeJZnbAHtMqLWgoLtodo9E9VSNVYnAUnqQkqRlkTB8r/s1C3I4lhK0o/gyt8JTL/+
YpcLk/S6XEX/Jh9mm5lLAmwn4TNDMy941yvKp4ciOnKwiGlQXZc3TOgNYWsOUdQ2V7l0gDNdhpVN
ljX5HjUoBZQWxunwgxTEkW9x/fAjwuYFsWlBSqYzT4T6Ox2B29aJFHwpTFE7nCmN4wQQSXYv/Z6J
GMSOq4knoxNxBNoVTrWZAV707HhdkYnBzm/sO3pS825KuphYl/1D4VkJEtalMyMmUXOSiOjz5YFq
V33GDSX5ajEHvUENtiRGWj9XilpUn1ugDsL5feuR3LfRKD0WhVKrN3iE3mQ6tKIbJbdeUaI1L0IQ
AcbtfKKxCHcOyPcZKz9bu98wxSztpj8aX8SlGN3m3ufDH5FnX1Xr3VlEuCJMDUC1tqG838OCwUYn
GszWrKt+YgwVmmL391ANPO0eXBmTabZHCphY0TJFHia8ufaV/cLc43uZEWosv94XdKmYmMu+p2dz
gh/lelFHc4JTth+yIt4yZejLosirEUcuMf2u78hFKzf3DKKpLGA5FmltD431rFU9HwQTByNgF/Nq
8b75BdbJvv04Fo0pavXinZH79AAwteafG08kpQ8mRiiIorZmhLMuwYEgLLIzox22VmihldKe04C7
HIAopY69z8Tf0Y6bt7DgiFAs9aTE/RzInq8LkJAKsdy6Ab9shao7b5Rm/2DX+kyfdS6zed4rrbj7
qMcExNMePrqVBRHXLP7hy3H3cZU4dgw7E9zcL5BU4gn5IyTFr3K10WeU9fjNVfwVe6tdkmiK/i6h
ePD7IgHF6Of/ryUmV2WZvXZr7KhMxfozvrUEcTri0CKkYbUHzTE4FK9UjSxgFgFoyMeZHUffhMK8
lllXO3wHoFqnheadwukIJaDYxQAxbWWgZfIXzkl41NHINq270FWcEuxjFPJWU4HSy9utWfUJpk7V
cNxppwxjog6a70x6QXEhk9Kq4EObZMwP6Al4X44GUaeyqkV+jok7au2AS05U6a5yQPUoedVKZnAW
Hj82oCzrMj27MmuLSBagC5Gse7T3ynOuCsjsWodlOipyxf4D3HwqMu9vYoIcnhD/Wqoi2i8jOAjN
S/vjq9vX2eBVA9sW1FetieqydTT3m5KwSKuxjjC8iNpNqK0gGXdIFMg/Au+w/nG0UuBUjfXJVxnt
OXgGTxYoLlWVVTbdi+bJQ56F+Vg11UlcBjRSqoBLB4prhrHVwg9x/YcrKE1RDSkbELbh2JXLuHfk
G84G9o2KE1x1PAOqsVb8Y84MFBx1tr9yBOa1pgv7+UzWRlR6yRULtvT3fm/HXTRbR1h+XDwbi3ws
6sPYRZaXC9vLROJzoYGCxneDIwNG+O42UHotzP8P4wGQ4nxxGCJjrvg7OIdG5v1wgLj1+4B2ZixI
ZfGe1KSPoXGkc3T0G6e1vreh/yyPz7BRha/Wq7rCb+unkQ80hoKGMk63VD4M5HKmGNNJgfP7JF0Q
zB1fdz44DMgtcujQYxfT6PJg0gAQoccDfNY/kn/j3ftpCXMsuDDemd6VjL9P+hFj/IfUBxEnMLMC
E/6e+QW4zyb8xIMROQy6dMduKJ/Yfe2zHF9pX6Sl4Vwb0b1se6yNae85R4T1jBuyVDxbSk0ZMRtA
F0IRtHy3gaZMb/mpdhL5taLBsPtQsp0C99gb7UtYWNL6zAcohuYBbhQIhoGI8aLn7GP+ohf0iklq
uwDg9DSu7Og8B8Ds4KX2E8UPiSGZ5ncVAL3qLubnRb7Dvcjp8ClrU1/NFNe82hnP7aP6jTaudrmn
22chqbPo394Z/ytwNCxchg3P4pqWVM6PQqCzNRTFMI5gYxIg5ITxryZag1Htt1d8n6iUOtxbSFSW
CHiNySsemG72fufyjfIXjqX/lef5sHyG0INieT+wSH1hEhclhop0R8j1spp3fR7skz+jDa+X85fW
kx45xrSTgyB0JE/2/CffUA3Vz4ahGQWBqGnuNQsnVWFpacxFlu+vN5c8WgMBjX2uC0DhShJMOSJz
ZHf1M1D5bbXx3D3rXkIMUKi7b2bbqHRzFhLHaznUZbqjXg5nGrJzDLX04lQjwLGtoNPRhkcr5VyD
qToRZOm4A2z8BXhtOrlDUIqBmctqh4Rtaj4RSQxUSB916NwiNKvpZjj8H/U3jleOeJggOWgPn1Yu
OYU4W9uyRCVgsNs5Tpm3iSMheabW3Pbs0OTJM6Ja3zHuCahLcA2A5u/09HYrzTnz5GpL1CaFgo6W
l3awpjZmSFddLzBcO8BFUCiwSbLhi5tdehRnGJ0nLV6Y2BhrkcVkX1SB+YtLAnNA8S1PkpKcgvx4
q8HMq24E0naAryovMsPmzASAQ/202zGGzNHCicMRirvZEWJeMpnWjVUbKxZ5Yz0u45MwZyEIWFcj
D9FgWpEzrmXiQmka1ZPbDVBpkUWyjiIyHu+ly2ypoWsD0U2hIS5OwdYQlYmJ3CLXNGaTqynV8C2U
20p6xSOEIU3pycLz+iLyL3r3jtwWFACQWQvYUHaKs6U+w821sjXHF7OOtNuXcN6F4WYKFQOK69/R
hXC5kDSIJRA3j4aaJktXbS3tatPZ8LhiFDypQ2ff+UOOC9Y/+sBDE9Kf5uTqzZNJxpULHX4k75tm
/eRnTC3ArjhRmsuBGW85EM0M3o5zcRxClQJOh2e5MHal1a6B9DlGpo6vEdxM7C3XVjG/2jXIDIeS
X/Bw5zjQ4KvoGrkTofT0PbM4OdV2QPOZEthYX6uzRwo/Dg1mLmhX4OQLEpdmYp+iSpsD/dVYN6Qi
20GGfycVezqeacaskLrEMQyH1KBiMEer2+FMlxm0U+xh/opzVwcM516WroLdWt+XV+Ei0q18HsrG
/e+5xeAqLMv9F34jvvoSAUjLRbQZAmy698dHphSbBV2DWnpvyiMXcs1/ZF4/N4H0k1IlThsvIHln
tvr8KeyBCMggWpsvcOnKWg+1C54RlIp0v+8Cs9LZlo5vfB4MHx+zp/C9z7bUzLr6/wk5nLaNZFHo
f5z9eHzi2sfI5qjNKu606hCD3It+u25XB9CTReymRNPNeJ6vs56YnlhicI4lytV0vaSAcuzGZhKC
C2DqLzEFoE9kouizaCkrRtqXnYnOJzsWxmq/qjQ9KDIPsfbXWlsDYqmzCLgT92xOvDHPfHMbmGje
4lf6JSyR4bn7cniPBBOKyQg5VNQ2dpzfhK5Ept51VeNnhPuNizHLPELwDdv3KI0Oo5oww47tySge
w5ctHMmRYoc5Dn0Cp7EfUOCFRUL4zD49LBDJSWu9tYJhVYNNKLh+Bj8hKtyrB7aGIrGKJ99T1Nf7
or+AmwsGDjbeT6wh/WSyaF77zitBiGQiZbqIg8XzqYYgzFywoOC6m+BKd9J6d13JdlT64gYSxPqq
cH7aXURJv37RuDt18o5OcrQYI7CAh/1c6R9U3er4nmwCQKaUk/qERlzqGVHGdqM3iSIgYNsmlx7W
nioAJQ7ymEXCQsk3WyoCuo4Ee3uo//568NV4be7a81patkSv+G5Dj0Uaounv4F4cecALZStwpYxE
t29XMMR3+HL8SqGNgVsIqY6osGSmiMwKpwLlqipI5OtSpsWMvgakdtg7l2BeYhadFHo6FhXmxK/a
ZxqqoIl38ju/fg0IXKNzzlOxtsz25AKxPYhM+xwn+6dIUVrferha+8aUB/klxgXl3XXHe8CeCNMV
qBdt6skNttCoBaZOsN0HvZ75+uDep00Tt7lYv6rABq3gxMz9kImmnqAMBdIY8Rlrca5/rczKNg3b
EqAAnkE8NjMtHPtpBCmETrD7NGgXkZO//xO0VlL2O1U5f1utvbSypkbmpJRpZMO18UziNDbbjIPY
cM6Qonvwa1tqhTMznLm85pQqi3gVVw11BQqqlAQ9WB8FfuwOfEGT0BQaaaCRRYn2941fzdJU1AQY
8yhvN5AMG9N4R6YpN4WV2qALB79Kz8/O21eHVQ7wPprlDlX9mdwPy58npszqNg+UWK/fyfyFGvKd
qw9ZTXPcSuWnM3zr+c3q5cBhfplGygkFgjH21gn0+adsPtnodko/908dtTlBMw5J6b5391RgoREl
Pdxp0byDA+29lGOBZuqf5XyNUoPcXr8rFDIeW3uN7LX8sGR6fNXwvzhj6syyhPFwrQBQ87Z61yFA
g+dGxBLFeK5GV03NZMByRhiWzWUp1Yts66eepj84B6lUlawZsD6yTzhL7q6jOMqnaahqCOzhpIxK
iqr4HlD6dBX6E4uYevzQ9qhVt1XbhVBDTuBlU8D/fYoozXp+8uZcp0sA/pK+XxYS+bZ3+CAftKv1
S0r4pnP+/bmdl38SQz+vrv70hHAvXg+rWiqBaDNgxLXrmC7SqVsGa7hUNjZlKuvgbfvnRd04WIeJ
jvHFxRnfbgKDmtgn9Dc4ETHKTYHt1Nc4CGe+KQGJ3hMNkGcvtI2qmQ0g4iGV+o0RgWzYwpYOD1W2
vAE4ukpdTEJhydBkXtHzXpfKo7sG6b6xiKqEczl+tWUj5dkTm5BPGDL3vB+CLpLXlYD50iCXFHks
zDbtn6dJYDrwBGvG2S9XWPO1b0Rsq86as/F2cWNplelN2PkTpfrS1VgPQbu3arGGztEyupibYZpf
QUkmu6MzTfZulo/UMKwaglKbgv4RF4J4hxHouAT+ZpefFzw2g3AoEP7o6dSXMmqwUTls6M2AZLaX
3CA7YD8tsRuZipg8VklRqMLLaLxLCjkL7V2Yjpi0RJ+x85EF+nkwTHmSVyf2qUS2ZKmSM0R3L1Zn
S0suH5mSCFxVNdLcIHcRFIyZJ1a9FRwG3CBLh/aXxXy2py71RpTnfOsj13SzTKNZokD3WhwqAs3J
0RQji75tLW682eon9hFfnD6QxK5G+LBoYV+mvJoQt5Yu2LE8ech55kG3SW3HJ16gQOuwNy5uj8Nf
5EjXcNYg2A+8MwOJfFPmyKZH7g23oDweRRFBhys4UjgnyXuGYcJOybImF5qUvFDd/kPvOHsz4vJU
Ng/y4EvBbNaIpiQANMgIBZqs8lpKQjD6+2hGS4ssunQuF7aOQXd4eK7JBKN1bMLaXJesGhn5Q4gO
ljni4iJzq/SDKRJBjwwtmOaeOszQp3OGDEeVu1UFkVZTaARR+dIu8lmGZZ9P6EIQ9QLZ0LTmlZor
1Wzl6mLmogCLqsIV6lNslQQG5sIW1H1BAkZ7XFbmdGCEewMi08tO4+UjG4e/S8vHWH2qI+e942sS
BvRwPx+F0+kGPYDUnjlRVrUwbN6p6lzC4Mou2867Cm1d1nsiGj4N1XXfiNh8G1ybPzEC6435YbvN
eKQ9f/50iXFDHaHyZGwF5QUogUlLeMyyAzy2xfKSQ+AzedI3wjGTM15pNFgo4xFdIL3TWQJCxu2x
XKK6SV75Ss+iwoXpSPvPZDa++hlUWwpMEYmEENtDPhzLCaLibtlPqlusiotCKDU3mpDvYivVRKQP
66Gii1NvR3imTD5nEFtSXvw1WCTp5fobhj30gHeENKcLcyDONPeD3wELc6+SI4usE6A8yC/kfLVz
E2ij8WNuLUZooLK5vCn9mf3WyP+z1DfEOozscGHJnRMpVOm3Z6tGccVpFNiLhImQjSavbcxyK+jF
BRmbhIrtjd+mPx4TTb5YxIUGkbDFQNMxFVUZwZIWqwGF5Qfo1vNpkhlH4etaTzhD6DooigKWfZEG
Uwt50km657tY78EEm5IVE+rUqC5tAiL/oKGXvHwl9E9iQG4CMoQKfsqRPN4W5yecK5srqxV/CODC
qm6PP4eQcI1ryOhc2g4Iq7+wttKG8DbOzb63ubl1pVIhKxMBlbNIXjwu7QUb5lVzYbGdk3ZsLJMq
XWyreuCgoE0dPPOaZbhgwKjtjCCp7DkSjXGg4ZyDyedvo+38BUOHcw317CgB/I4C1ma6DhulkRKh
Ps1LR+ZTcXQxKIR6jPix0YHosDeOcrMSXMwrMs8rvlHzCumIQnkCSGnnkwBIG6cUmxLHqoiDJcgz
lTchgmpHwN5HKaI+5AggFeZqHGjJt4FybSTXLdLEIQGC00aQg5bfNt3JdkwJZnaimS82wnfajPzi
QnqFQ9ocQWQ8E9mMVqzzX3W4RDM9zDEbdBcSyuaAlU+KtoBhGW6ugi4OXNwWKXGwlkoG19wUTcyY
kAOZRoxi2/b+zhbpF2szivq4bpmVD9Ga9LQ2gjAQSXYR7bcS7em/eGV+HTUbvQgDy43XPekio8YY
WLYxKmU1/PqGmy8dkPaEKIgGT34A643lxMnYHmeY9GW8PxHuROr7HiE3KzOkyarjHgaAAZ0BxTbQ
bcG22SxH5sTeaMpFs1iT3tEdbN66BVhfZZON9Il/Oyqad+iIp9qDTF1eiZS2xAsegXbnsu0+l7uc
GMAKIYxpzxXK8/nrzBCj8+XM4lVRUXpbqUqmPVTaiamdjHZiE09LRWKrX7vvMJ1LfzFmT+i+OCzd
BGSx6dQyFVkyjmA5QBoaBI1G1fE7HGrEKj0KwnvkYBP9YnLXNYtommDgeV+3aoK0af4Go/gYJVg0
p+aSqlQv2AzKQhsssYmztIDZa3bKl1NFd4oL5h9u5qisWjeOU+ZZAaagpSdso9aMVUtIrIZD+owi
pGndyT0SBKSQUSUCVkpu9o4vn42v482MEOrg00Wwy6uKird4k994LSB5KDiEVkWV9bcvVx0AcHOK
sPN+rv6gdJbyjXeGZuk3fg610wfSkKsy18LymM51exntXoUsbgBPEq1RPH7JvjniAVoLBXyZRoDI
8/4zDZerU9zJOyPXWuxP+ej1ClkjHpNd/+1TMBD9QhA8wigwuH8+hWNprFQi3HKIeTSF5tfC7Afb
HwFEWdgNmdGZpP0GN56ToS5tvC97svXgB3oSyGFrGkx1TWOws4/UI7itEHUgKdFsjSDXQ8j8nGpl
QGTEoUcn6QuUwnbgZAkylCPK9mL3PDtPOD6vtZ1ABxSxX8Ph7XSpH+FYS4tFiVX+9xUYlYhEJIyP
tLZgAEYQ3ZttvTafGMwWyznpIlJRLY71BUvjdFrT8Y0bqUx2MtcNM679MCqhVXXXj7z68+jbzL/b
ur7wBkNc77whfXWGXwfY4ZONUrryFnKZIZzvEM+iZWSOngVE2eYqsR0k9PcLOnqgOYpee8QxI/kk
tBd3vy9AjhpnCA5bdXGX2YXfT6ohZRGQ5jgBS4x1TGHdcGveUj3NMHdtdzH3Lp/QW0E6H21kNZ8+
kqb1Otm8I2KUJrSeNFEVUBGKdaJesJLdtIk8XpoD9Ovf1mPvzzZwIQ9+iduW3VoLbb8e1nhWOaYK
SQgI52R5GsvyCCkk0HOV8YbhaJSFfKtsL7VaIR8UkmNqlR9hBqi1+4TlW/XjplsxITcxr4lX1+ja
6LELd3QM0h+QhZWj0Zk/wytUCJtHGtt2VXxAnrQFwnEY7G7Jnqx8X62vDwW2h89APUHc22EJFvic
10wXYwEIn8uWejoLKf1CxhnygARsYsKBAIiNSkugekpsbHCnvs2G/sSvRMEYL1pln1zvWUNrn/E2
+zFT3sGA53NtCe8VPcL0PTA3uUQd01eJF0xBJ0+7rqpNPVls2o8ypntGAtOy3Nie4Dk0EIvXFHHO
x/NN7nQxglEpIweS43kRbD4JpKt+xrosEXUGclNz4Obz1fB/Do5tv8Otg57RwonCgWfxjd3m/3bX
Glq+b2wRaPiQDzakGOnG+9rDnZ/U4kQmHegnJYbIF/nel1lO/ODL+S4c+aH011/rWDNsN1oXzjWC
db0XjxVyW7jAUhOYS6BY+fExTwJp9eW4xJfk7BUx9n9s6ePEhwo11dDtILZpvqvX0qm1Qzwnh4pH
eXmoiWeorP8Tka9ZBRkX1Vfd7q1LQc1cTQh43ZsML5A4hHw1ERywyIcQUyVL732UoPp4CCiqE0Jq
z4k96torfdGJ7RgjdXD5YMbHCRoCMAGJmq0po+sDVASyuXfaRL4akwC4qmN9urrJ+awosEoL+5p7
0TcdTGDCfGF3mQHe9t4X8kD7n55ezFDRtmLU30p6W9BV0bNwFsyONoJwYEQGYvVFH7k00nPzPTkp
Vl/xkqS/bLJQJc/vieMtY5jE0LGZOCEBr/dfbFkhK9tIepOUqhvDP6voKMTflH1m9eeymKUVBT7O
bCY/4SGDLqW6YGmtZYCiyIgIxBy1aLtaCwRiS6qTGwC7RROTWKe6i+rFzBCwN/NjdLIs9/enZF+e
eSYhxLwfZvJQx4xh4V4C/Dh4EPbneM/2dCAxxW5HWcOG/VCxvpXhPoYguE2JMaGm9FalZZ5XUZRb
kBB33KgziSKei10Adqeb9+VlZKdDI4/Yjg8sSp/U3JW9E41s1BVfqOnWfACePg0wpgAnGoPGbBv6
NQfI2a8N1pver0pTe+Waw0qiFAtBlTsv5tSyVXo3S7npkP4h6k6rOUpMdBZDyq5DssEVnMb2WH/j
pjFwWArYXeksX6PE2YWkOitdHyzYQngs8yyESgvmwjNFzAAJc52AbwIcVBfFyjkkbLjUgffiGPVf
EnLU1ZgJaMfL2iD8rZsiDcyg1CQEY2aFkjboWGfnOTezdX92KhGbXNxUGmQ52SjTen3jCit2mdXf
QwqLAwMdNwvlSf8Ba0WpOWXZwc7Twr75roBbolfTJfB1MmbG0OIS8KrK+CgeViURfwRnUBUkg2dL
rtyYUuLz+hP1gkZnEAgUiz5BB4sJcbePjqekYecPAdiem6Fb3IrIOaLg00x/dHPpCussSb+IiVVc
jIdsw+qO5bLJX0cJi8pssNHYFsaTIOalqr70rAOUXMGv4ZQ0AsAP7uBsv4yvLP3B8/XjlFbL+qIa
MZi6JJKRaQ3xL9hkHWfLW7NuwwWXGUqEx0/3GHvED2xiy9XF+N0+oFy7h2j6fMRUzuCiNhdnAiSh
C5Dgl2u02a+F2w38dTVwP8TBqaHHE9L2geLn2kEEW3vD/1mbVA0OfB2ZLr8ne6NTQsRt+cDbCRfH
I7HAwv4GPR2VxcpYvaQyx2etlI6B6r5V6Jc7scVBbMlw8yFDfaZ9zSI+ri0Jy3F2pSBmb1GYCdLp
eWXMAnw6+MzfG+uri9l8CVMiCaybErTJfwhCwqliZaQ/bGnjkPkpY9VT8Qzbh8bilz/1fsqmm2Rf
hnU6MiTE8fzCMk9NZrthEp2GiUtLqwN5nv8O5kPnAJEAjq4pWTeaNjPWG5RWmp6Qt8Lx8eadzQid
TaI4ur3Iwx3F3RPENOiEAzX1dRnNQQn5jqJrHKQD2r/Zridtol5DmFK2ATw1XusIAfppUmtq8vQr
U/Qcq1G0maSgWoq1XdMXfvxpzRI10fR5ezKc7qrXYRarhfIs/9IAkPJvQK5558E+dOv6Ys8n+ago
qyxfrS+AjuSmnKwqamNLfgmWjWNPT7j85LXU+qHWFDgIf97+hPoYyVLPETxqUdBrGwg4Y2TxKUIC
6efPfj5olg2Y5ZZrvICgq/hLtMVNNKTPtK1OUzOITg+h1/KWpk9Nup+4dQFPYdMBxENAoe4aeGYJ
vTdhtGxb+M0Ujxa0DsJ3hc5UrNKqaXIKWdgooiJo4D0k84an8x747AWIWk9aMEz03p0lJv6S2PX1
Uyf9GD2zvO3jIJAkzhaikDegjMOyvR+niBgvfIPE1LE7aAx+8quSxxZ9ml7y95JGXsCiYNZhLcF3
BjAHhrbtPVYEGrVAiqrvcxFteK9exiYSroewawHEuBWceZj+FnkbNh91FWAuZENWRuu165N8NDMH
a1fN0ZAgQunPBmRe4hScMt7/2HTE/s7TYTAJgLqB7mocYBNP25Rub3gxKz3rqgaXQeIigTdaCFuj
Ypw2RV38NLIsOwUKlukXlw4e2vdDg0ODEsNggxD1J9zjCnUiDXobm134G4MeuNM/OKzyt7xDL/Ew
BiO5HouCIHafopTDj90n0JaUTjl1cu4VmmJuXvdB15b3Vi4Zfmw/zNoVr/uqTIBz0mm2xvCDbueR
+iZvJ6+hwxEDTUNIs128t2Z9v9VC6w7+IX6gk4VUXsZTsAmjxLgWt69R1Kotf5kvhrndbnxTLZ2O
9eGprDqNyO9NejAfvcxwtYaafIEKL+O7+XJ3C+DfGhh+GUCmW51WBXQwJ1WBOxcReEQiQWLRxUT0
RaHQ/kiGBo9J3PJTTzoSghK04PlChJSOnWW7VqvBKLw2SsWQvDKOEMHHkGv+0vsFOgcl1M59ZyRw
rvgd2TL9r9r8gENvcBBA8R2NNT2htO11jfSAsccadpsmkUizN8OKdBjCMKNQBqIxcq2w/Woavudn
l0kD5DCMx7GQI1ZZ76+Q2GhmV0vU+/8NPcwIPa8r5JXyxm++6q5EOXZAFsEfPodzc4t/h+A3Q3Ln
RULihor1cPqe/AkNB/kiuuMWneCclVjNthm+JXK8BlScX+j3N8jKbhjY3nQTshidqFze7cZo6tlR
z0iFIwaWPKolCWjYVyoyCcccp4eYsTpX38bLkzBoJ5xtSpKZnNU/a5DVMHWAPDvZc3+p7Etf+76S
+XEP72dQHLGaZXZSmvCyGScrRYXPrASVtP1S4g6DAwLB1IEb3WkKNXXh5lnyAAJDi8KJNhSaBa2r
DXZEPcFDyONF6pY05IZOi4odnnovpkOXh9662Nnx/nWZTvni04Jx7kDvBn15HHGykzWlNrXqGAKb
00hybZa3D19gsa1ds/fTwEzeLvJOPrKPIn2+vMUcXBkqvSjpU9VzpR1ZAmC8H+k+iSAFdQRtYavH
QUR8bq1RY7DrzswT9Vievmqg0fRVAqMITG6akhkSbJx2/1R/FMSHK/z5Iyjj3PfG/2pEEwx9aVA8
zF6SQ47WPtPNSB4aROMXMnlrkK1HIVUKyEbXutu8ayxVRICx78ej1FIsC4ykMCwKWUrZIWEI4OKY
4Dzunp/Yb6e1paVK/8WvJRcYC5nyg1ta37pF/VhpoA0SJEpdLk+9m9qQ27tIPwYrBSTCLANLciyn
uq0+n764B3UA8oX54lMmfOfwwr9T7vraGe0jhaHUlK/JWOFFv0/Y5dcZ6vHnODAjSrrMnaxN7NkG
DUw+uqrK7QYOPo948apVAIe6tgWAC0+4Oe44SO+dUVXVBAI7qRqALiIixq9w9YYP6xJ72m+9dYSe
P/HzktrMzLgCGQ9VasColV+0eZoVvpaSErFz5OPcOTwdzaAnLnWlEtW5nfGUDZwOU2uh8fibAoIR
u/VGCS7vFpZtVuflpxe42B2m8A1xv5iPKQX6PGoEpjGd31ncP8yFNVzdszL+3n3S37TdH54bvOlk
ecwaRdjB5RsqibpP0qCy+Meye3oqHWWL18rYu4FQEv8nAWGGOR4MXs5/8mYtnsHj8nA4vIoO2l2h
as2BA8vBpjAHefG8nwwi+QUZXwX3KmA+vmH1t+PvUcJoIShI/2p01+8+yFqY4KkHrD4sLDfRbkyR
nseyH1OOw58riDpLLgBH9G1FEbKJ/K7bZQgXxzEDQLaSmfI+t4OXhy6hpxeOfx1AjQDGQ5V5Kob+
E1OIfH8vUuCzIyFWxl4C6oe2WXwiSe1hfYSXjkIZxvLTAuMSOGh+PccoXNgaDf4PRauDzaC7t+5V
OryZAmqZ4odRHvQbkrv6xThJXe4lv8OsSOy3iChbI+lA+GTQfuIM2S4YlasIceBQkBP98wjSK3ti
Gh5IhKkWjwdimaaej1kxpmy1qYLmwQhgeeUpBuZoeEAC0Ubu20joWm4gpx03T0dvBcyhwkz8lIo6
JeNOZSOrAE6zXqRZYza2hfkl53eDy/nsImPVbS/SKtcT69c6umD9QHnlLANK3Wvs1vu40Lx9Gugr
LTCJdLPTfjdz/Y3zC1rvLay1AIQ+UMz9mH53CqSLcCuiXnvi8XtxNsi7yIN8uz6y5q1r5NTJXaNk
AuztxK7VwGm1c5CUGCgu0CfOEkuZPxiTXT/ReBBzZzqL7OlfGu3tqn5dvMTEAFS0kXhZuAA7TeHr
erbgz/n5IzHUPd0ykWPDbjKkaMMpp5TZhny0pngZl/Z8zGx3MwjK1S7LF8HusGcngG9px0o4xLYH
p2yRQ3REw+N0uWFtP3svFu0eGayoy9MeihjAvScBcJAt5PM6RAnBp0DwayiDbWwXIiJpL3taX4bN
JL1/BfhM2pnFhqo5E4wTnPHX605pEyKRhnr19bz4y/GIB9VI7S8njOjbL1wEa8XN9hJFZoRwZSfi
yFek067sofG6QkK/FTOWu5WY8Ff6qussowmiNGtoqdvxRBMzBHsRWr1rjT0eYz3M57j7BpRf+kY7
GWcVHiR0iZdcedYaLaPT9jFM/SJID7jc3Xfo48t/f0skkkr1TCKjIqoi7V1vSUNiXEGGoEv/7Z5t
9sqCGNhOfIB+i+oj/QGDYqHDskpeygjU7hLujLyzSQuYRxkDEsSVa5AQH3sDHZ5ESdAnRvj+egGg
frpqs82fj8Z+ir8JA2EdJS67rnMGhbCczzrYAg6iz1STZ7mouZqUWIrA4bIrafC/Fcj8cUDncPrS
fVC8Cv2YX7Fvg49MDyf2+8dZ7rYX5D9k8ClGGnUryn87CG4UJrfpjPf1DSS/DdZXbCBaXAFwH49J
5CQwVPKWWEmi04CAWUAYtXZtFneqnwW9Ua/DjIqZ0643WCi6WaN9KjhC+PeRhEUdFreKAXgqf5dQ
mRQ0nMdLp1ves6SfICu1t4bw5jSzQiM7Ulh2Gus50RPfrqjCDqzlYHvKRlHHgu1fDN21ZYsiNBUR
uGNdOsl3WAvhOsTNZNiTVFUnLTUBlIboBs/uySThNev/WrqeL/vYoROYGSeyOdXnwh09IiK+LkWB
6FZHXbwPDQD7g+Pss6RPMfiMTv4o3Z5qyhAzfIzTsZCCUU2iF3ZRMXHarT0DiDylvNXV3A/04viC
QJwRRV+mk7VTJHzDuXnkX0VJVljH0YcLeOwhmSNqWhGfroBOlfwyaYK2fUXX3H5m1CHOSCES2Lhb
yeAi6le4RJd3+qSH2AveC6KL6Z/ILy0/YoN7JqPIKWitsEOJ3SoTBVytWik/8PIMmnvT9nt6CVS1
7duyDqaxvZkkn+SYfz3/PxER9dKcKGnCnQx++6hyhd2HTg03Im+kiR36iMT2hAIYsNyuKxQlGXcA
T/ZlHe2Wapa0tG6CS+cLeN9uLOYEBj0/9YYV+0Cir3dBVqokzs2jAsB9GbnFalsUM3YIyMS1VJJ2
qBmEtxaEnT07R+p6W7vpYJhvTTg9ymYbtHPjg8z38RzTq0JXlU7j7V5z7/t8d3YACmrJiS6QNnbl
L0oWe2XR4OWytk+9musIAk0V9P85YGKGNBmWPShTHs/7ssPVqOAlTyWhgVsF2Ouuzq+PXQGHWsCW
bmIEf78/tRRlhXZskL8u9TmZkenlGMIYV3WPvW5EXkaCYQ773D3lAtVFHs7OopmWnsRNK/P0vLZv
QNhNPRUZFkXodrr6EnjsaXgDBcAzBOY9cgYDlVsG9PBog34Hs6WUH+fqrTjVl9GmguZPdC1raARB
cZ/hBkcN55YjiLqsrVWzraO9rTVJWaUkDrnuKYpye85uHvYEbLoRvsRNc/yerlPXbR5KGEo6hfin
b7XM3EPAdRNLjCXNG65jvmGEgeoiKx4wrlsn8s4ORofaadvqcmdxuaSqHmVn6rfERYH5exUgbKvi
mYjdl62gmeipiMTSqpaWJqxe+pdvcgncUXN1iQZ4Oq6mO2O+a2EvSw0YPFZ/Ikz8PqqeQ58aWlyR
a5cHR4ycQqB/vc0JtaVWYzLdXkdyUhazLpC4dPtbTvA8oVgbKZuYRUOLaLDjY7SlvXx545vjvEDb
6i79unsyYyVglAR5VvcwoeRpv+ad+NptAbNCXbvh89jTDA2b/t3muhzx0Fq/uPYNMv29vuAZc0aw
Iv3z4nNETHaRXHa7+1TNbxGY/dtBjEMFKR3suJxNArdVbTieShk6pWRoZeAekabj7KohYgEO2/dN
faRlhCnYOO0VEBd8QXy3soxvpILyvD4s/UiR0/80y6sQK06EC8Za+QENqFo8zAXezReCai/mqXCC
vhH0Mpwrbj/TLcJFL3s10NTYdkmp5v2oH7mXguWnCnQzFaRm8ePJUZkY1ID+SPMoTC53ZQwAjER+
79Nh8czVV1xo5Rv62LtRiXcU10dvhZFu6YOVjeO55yfCvGz+kH4+sWjPeetKI8DxL0i+yMTl87oD
G/4C139CXkVWygyTw1AaY9g7W4fVTbdGUvVTCq1FRgUIWENS1eXG6yTTyJKU1+mhupuHRA+oJWNE
48hIz0EI+v1IAbt2wln8fCbif6X2kwmE393F1U2pfyKQWrBUSOgdVmHxa1GJsTQ+q20XRhBQdeQH
Po+/YMRIspeI+EUWSm5FUkDvAXzFY7r7MAG2uAtAW4BVdlWLTCfGAeLYXNkf4KuPT/+rNspzAzwo
EhJDw2PMvkCekzDTg13ovD/kS6/zuUDX7cPq2FqayqFtFiBS2yvsT41hpADxDWdqyAhJlJMeMNR6
9vuC1k0R0I/q+wFnz3K8tyasI6EWhFkPlAkVSOQgzFMPwkMsxjxkwiiskBnrz1rsHcHw94mtzL88
SF1amTIyD9S57revjqV4pJf0LpgfYWieD4Kz1jbZwg64cpRN1XPTcNepFTm95Q//HSN9Zk/kiIJL
ksjGxGICplPHh/RyaKY+ouEjds5JCalUpW6266f8BW6tfbg82HGeC/358SILyJ8E3KFQ02Fjl9zu
V4H0Ktd202c7uDEJsJt+/7Utv5Y/E4uRYwVh4/h+fbGmvfpqKB630LZNn75LpS0UhnlVM1Oh2AVC
0zQcQepLMH68+VhBVGGiIHdFJ05LYq1RfcRc535OI8TDwnhxv0dUYScg2zqCVy26HRV7ALsajNYw
zk1VdIi9oYwuStihw1bcajdqxHZbjDZMN3Cjz1bn+yGCw5oB05aWFnCH/z5BWHLY8CBhwMAnw7GG
/hs0rWJHL3Og/l66qxRUVbn2yx9V2fDDYnmQRSlILOT2PdpLPv3gNXDQTCknfG5eZRpdtB3q7qvV
biaDtL/QHiENAiylwhA3IRNpTImcKJGUniPsZMzauIY8qhqhlBiQz+PQLa9h2Ec6FMfq0avSQ5ei
hsP0vKeDX4FCNX+H5CqUNQqujyMWJsbR36IoPnFgls+kCda4AC/GU92Zhs2jG9+x7o5uZxPynvp5
3yW7UVAXVAAmSp/CTkOC9u/uDfMzTOG7dhhecbj1DDzf9V4ot6FG6/sauvDvNKlDTSiW3qmHeX4J
fKMS0lT53CSAFv9OHsQOVJjRo9BeA03vJGAzUinF66UhUm2b/YLRbHsMvlrLD8bDWHQsQk4z89yI
q6eGyNGWzSAo8WOX1axg7OF5XEJHupgS7TfqrpY+HqFT34smEWfuCRKL+45Ep5i9PtYEFL8s9G6H
JBdi5IiIEkQsNP2bhcroq+C7CAG34u/EggQhlUJPPa449SUDXA8htsorKHTybwzDBBS9hNM/5yRo
KoHPzKEUAvzeBv2+ZyGAwJMvRE73987E7Abb/oBlwjXZqVugsRf7iYpfbzyMxN+bDpkrthbJyhC9
nccEbTBS1T8c52XZQxk+gkmUx7/v7JnESADBm7gH8T1dvDhhrK3OLjOmYAqlnV4jJlOouBZE1XKE
oMF1K2vfKy5/PXQ6CnbcBoz+LE8JFSKDFkbQ5UenTMhdL0Dneq5nFOmHi3da50BVypJ0cZPRNi7z
d/Ac8UAyUWkwjROLdN1IsRJUKVyNwOhblJN2zlsQzZ0KCSgOY/0wqzJ7xMUx9A6OJoh6j8ocyGgc
wcmG2g+qXxaPHEV/FxQMV6FROrVzl64t/m7oB5bUTMn+B3Tr+XmyEoc=
`protect end_protected
