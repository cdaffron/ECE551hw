`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U3k7g85HBJ4qWkgpO7ul7j4ufWKx6HNC4WMbbA9wy1W4jHLeN3ykMzYx47fIahtvBfmiQnKGuxbY
iEqCQIOgUg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ijGZJW6yWIJgkmaQqBdGrDUtEfIx64pjZL0ZnZkmop1EA/6IoeHHEBTiyU4/h4z0fEcBdjZEWrhZ
f2zusR0KKdOe2F7rVmNvQy1YyRxQ3MLzd5fOjJwY+amKNcx+bESq+LoobLM+a4YGz2OZvdmhx1py
ph9dxG+mJsxYdQ0gq0c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lwGmhC27U5Vdd21KkGTmLGY8iaKBQTKwjm1pYpSRYcTIet59m10+/ymyC76YOztlun8d3MU0eF56
w60iL85D6DLWf0u5FEaXKx2hrlPcLv0BDTMmt9uL7H6IJX04FAdOSvG7mb2BRDVqadWv+8ZbGPuE
a9Nh66wDGCDiRp/PmLLe3dbJj/nIXWA4vaLfu1P05/0rd+vT0zgUSOuLW5szkzoNqz6t14FqESV5
IsrxPJgOfoUXeqhu8eqg7y96gzavBeDZscvEPdr7weqLSSHQxVYUNRDPG6liMuX6beR2QE7l4g4b
VNrJMsxSh73K/9mOwtE9CoJ57k/gRLVuCtOorA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RbEB8lR6CZZUV25zKLxyDHDPJ3DsGRXCA90gjYrjsBaRq1zdA9GAJxIIgNFWrGfjon3jPDrj/s9q
xlAlDMmTxwwCkUIEuwzl87x/OLDR+Fj2DCMQbdqCdwXkCvzH7OhAIHSwS+wh7fltg3j+sz7v90if
KaWCWl33oSPodUond2k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ft4wS9f+REJsVkIEHG7YqcuhrjEPj5a8oUsetQ8NhlENCeB3nV1ERswzt+UVexQPJr4yv9X+x4EQ
ytEwSdKe8MIxW/81+pBhFVCzKS+AamAQc0fQgaqa/2EYDKCgEm4SBdnloyeXra5RKdgcJu6JQH+R
q0LnOG3Rxtq4BEJJ88uhKUUHkbuUly9srftnrWXx9yYWv8b9Bgl0pn7tqm9YJmY9Kmc+dt/Nd9Pv
2AZ1VcUw5jxmHisdYjQjsBjpuRf5F/SxwJd+8d7vFyE//oFM1qgwg8D+q6ZskXaSOfAQEYMxtpOM
YrKC9mf4+4xshRAWW4fIk0zrPGibbNl7Jz9Wcw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5568)
`protect data_block
Epal8Ge+h1O7QemD7uQn5+to29d6JFGwc6x9m5j3BEK7CVzmkVoaaOJRItc0LP7a7qt5Etfmgv8d
zelodan4PhVsiWdweH+fvPNGcI3o3pituwtzNa5bAexS0guHHR/1m2DxnHgJ7Lxe1mvLztbKVJsJ
tSepqpBZh2JXGZFLztcq37LfvDzjKlTYbHyKP7+1XYeDBkNZr45mLAqblcdzZ0WVqIDsQXqhfkbb
jsZK+VqED0eVmhbQv2YlpGKKPiy1t2KyVDDFzbO6hnhhdYLcWsWhwfEE+2baswrOoWIH6T6BXIAJ
CKa6ZYx31NshvdnT31P5KeHWTkRGL6eTIJaI28VQ0N+ihq8aF6wqM1akyrAGuOP0au7uinWsPcJB
h9Uz8wVSGRHXAHOs+xjiWe6RxRzMXQCPOgwGYzZStuxBBoI87ZtriK7S9abFsESCiMQCU1FtGXKh
qw4TIwS8rHcfxFJQznRMDlGtOQygD1DgNMlI4qXzLUjWzgCFUOZg+AhpB3EJ+HTilYwwkakhe7HU
cayDDSGSZ8lqd9pebtkhDrk3+9i8It0Y8ZTGe3vMIq9DaDD5sk/iVqEQTitadUB5BFgp3B3qDwRG
BmryN9sbp/4PTU/GxEfTMPzv5mCeMmChE9+HinUOU2YuQstj4NBz4HO/X4ATJMqEFL8T/Wy+dO3P
C5nZATkyc/ob32GwBFy3P5OsspoghJp451ipwGn3aIq3MWMT0Coc4if2flUHFzEFkeEpHKK+0eGy
/ls0gdmdQhEMIZqYLv9ITksOin9DCh5xjUVfJXfS2noiqrHRXvt8+abJD8bVuKHHmyk0gB9L3AZ1
Dk5FwpqJgNDOTfKQvfMEeSUBBt2EkWnSL1DBv99ID6F0OYwsyhKxeDXNuw5TCgkTp19z2cT+X4fG
q7JM+eSqG1VZgok8tkNSh1uRIiEP3mJoc0aoonRvvpdCmEtEx4fYIYJoNYfhh6OIUQM7HjAO677T
3fqDUkDtJakNz3zVbjd9rujXKVTf6gxifUS+09Tt/jnAghXvDfGgBtQWl8QgA8nSpA2V1IrIIBPj
ewva+VsyhtL6CpOlcQFfCB+KyHPTh12lt31UuvdMkLkw5cmry75ru0xFbcsWNRLZWc01bykoMFuA
Xmp585xDLEe4qwQ3p7R7fX91TPwX9/kTceQ28giNzmvMuIMPddWtSaYnjTK0Ik6qhbfD7je20Svl
eRgM3bxL87r3Ny5a+IixMOf+bgwlBgqwSpUtbrIwVo+pbta0xJxg22+xsUyLqb8KxPYeuZOtOfVL
YNwghWa0W8zQ1Hp9a4pYswwyW858PvMfL/sgAz+hqHS+4GPiec7zfndSb99xHkTPg0+WXTwNBYoG
Z6wpt4Unmhv//ufuzr3e5meH8SEktnCAUbParrB/ncR7ipb7KOw9O/LGKRXQfNuElZlg+rCsOnax
3moOwHN3E+DUecCc94dJA85lGD1FNWtCKZv3Rua0DVvBAm+V82GXdJ49yOd69ApucuY/sLOggISp
JrfjIDupghKT0Qm4l0MqOzGoMkTweqqAi32RYZKyfR5CXS5uaLXzT+XIYV/nnahZV5t1b+PUE0Cr
CdjjbJLAmqGfViEPYK/9hdITwnaEnF6nBM35BOfvOCV8K87/BWmbcGvkBpSY04B/UFrqXKoLEWhZ
KRIJ8lNbFvBYZiEvXICsLh+BfNb9tc+BiXr0VMZhXrO47zzuPf6cB0sQRKadFD7FTSKGfiv09nww
HsGjvo8yrZZvp1GkIw3AAkdrFNdhOzqG4MGXOVIy1rj6kufbQSvpBxUmF9cjEzXUNudzIfMvnBf6
2Xh+5zRSyVk+2/HqPRb5XmEvThfoY18Vlt2O7aVkzM4vnf0x77pNI2P4STNKjpUqSo54POuXgrcP
tvLRYc3ylkA+7NUz000lebut8QSQh592J2XIJtJRW0w/vW7+gr8ayGolTPxfCrgjV1j4DJRpQTok
IXyXe8IYKl0qxoGIS5OQ5R+09fHhbZg7+JmXGdou+Anrw81tYCsI3edteNHmUSi8bYwyDf6zW9w8
Y4icVolhrhnpOmjOP4tcWENTzrY35PcJGCTowjT2sNBCfnxUMIpYRmT58bHnYQoFl63ckYnbCxmJ
vUydarrC5km2Zk44ts3ZwCX1iQJpWfXfjc1BpNYe8kao9LIhXS10Py27ktOSB6cCvfdfpe9Ioe3B
L8u2kvHMMttFiwPRu6ZkFTwQgE3g+oDp17XeyflDUBO9bvU7eaWveayLsTtpkLbQ9qWibYiM7piY
Wk/tJ/yL6kdJPHXM625rgXt0hnbmNGbIV99jZuJNCM4glAsujYtnjSpoD0MCj6L9c/e+mxxQPoxS
CMmLp3FbXAgW9E8A2cSLWRcZlH3Tvt237wwlsGuEHo/UFF7zPYRdFRlD5PtbJJGSlGDiqmksTtpz
jFusWqjC4C7UTfeGgszlU5OHTltVnYTsga9S7T/NCesOs/CNBxp+KZeDKeLE/hLEdO5aJauQw/55
5DpKRm1xo15eVjPmbfTD8zXuf0VVTfNrpo/ksQtgPuE7SGP0Foe0qxFDU1lCbm/ydgUxOGqZNoyi
SayvlH6cuXkl9eU2js7UbCZHaPPYxEkqLeb/xybyRSGlJaLLbqN5KmzV4ie1Y4YQCbITu6YS7zQx
W6hDRCs9fqbZ1if2HPRdUnubUMavzQHa4Of5+Nt5f21+g+2Vp9UqAIDyzjK1TOeSLBYkiUP6WRnH
JFQ0eLvfQEmxsTJjtVXbo1vRTUTR0frvEz0/RR9x+EwUdy2okFlQv36O5lf+FbUkV524lXzxumId
fOiA8AigsCbRZA5KPnbll6Fk5GN9J4IHMjdmVzfhmzZwSjzl8nF0R9c3zKrubg4K3tpdAcd0PYat
7zaMcXDViXOzskGzYBZLYy3FgxpGW7irWARca7tNOP7OWnlnt2EbRqyJwSr8jEgnMk3zMvroWrlX
+2FcQWQRWhGBOM8bHIAn6Y918iBCaV5NLXkiQplTy3GDT48+hA62+5HRr9Fgdz2CVTNDHHz6BVnX
whmmwkVC1tJnR9o6FMNBStECnF6PmutRaz7dgao0HeJuF7pX6fI+wkUAbGGz8bp3ZgOoCjb3Bbsv
rjzBObx7l62nTPba/jV3BmxxBPZpXvNFl3w6EEF82WMunAfz+9hbGwgybKO3O7D853dI8KOHOs4T
lwxWYIIfsJhisBXvuCwQ5ej6Tgvsx1TNCc9XiAcuO9xWBBdQWPWxSk7tqJVBA8Q7vbDhw+lhzIc2
92qfMKEcebe/rAFMhViTLaVF2i6zpiTjaANYXvFiMeUFkRePedOqT3P2dxFXTtob6wvyeftoBo1g
v/RQoin1iBmUXlu3SaOoCEoM8grhFst6hlrTMwWqnpqj5PFkZV0RpamcFrJ0DdPHuy4ioVWJ9rg7
3XehptGHefEDxIJ3u+oHaQpsPpT03N9azsByuyYfwDIXbFyQQK0Km9YcprbYkQXgH+vQ8GydfNvg
rj+i++FuWtZQhrPrp16tABBYiHVMvuE+LWm+0hpXpZhU5GuctmOwexNVVnpLfJgGD9dV6AAHOKbe
I25asD9Bvaw8PmvdAJf1IimoymyGa3TBp77A4phNf/sNeqPWXvvD2yQvkR3XBmTpp25brSNrdoCP
jVpBoZRRfdwb6cqndpEZvErup5D+4Bd8xiuTsrteIA77+Gf2HBno1GHJVX30rJnWArO76gMIl4ZW
0Cy7g+rlWpox7z6iaPpH+LiYWtUBFQGlOFZ3RUrxcdiLC1HC9PdHa/ctYxCbv1r9K6CWgVOBI0o4
htB70D4pRIYgVJhl3KtYIpifibUiPeBxyHP/um2hU6Pf8FZQL+51Z0n9vEcLB9CsTaitOfcmJStU
V+ZQQFyJQ7IWJTLWw3qsyJHkzaNmgrNBZhyhpHCZ8xDvN6HbIaHMx0WpuHleA0dbLYe6fp2zyrXo
xOvKlUIxveO1XIUaumR6VCmpjkXHku30HGE5dthfiyJkEmhiHULKgQPuKSBeH7dp4gLJkfVXYxL8
1VrWM6/QsGUkW25o5oVDh5K2Vs3n/PS7s4yJ5B2Uu/uS5dXcf8MCvltHF4om0Hzv2oVjm2KUQdSM
0FCfzmMz6hs06tPMhV6zTFmEozx9sUpPVW/2vmQRVs6aOGS2aJamJyYrfE5YonzOBjpzoFrZGBE7
aaoG4fQb287ftV7xhCsUN+VM+bCyXEg7SMtdlGURpzsPckS+GCtbajdHUJHBz1SiVlzgfgkMxvAL
0uRPYfHTMHtBkbm7D27nkJeKMN5NS0pz1YBfmdgWLcA+riqvErT1F28f+GD/+1DmgW8qlgkNEJPg
yt6hHGrSB7S+7JDBAQVpNdX7hmWMIA0E0iEwlqIZHNwJ9P7HPtNRqb/Wu8s3xvey7Lw3opEy1s21
TQIQLFIMN0MsAQwNhiAA7trYWZgWkS/AX/lJugiAIDpj0EeCZfh6XSFedY/ZyIiKmb74r2KRePhF
yBuMOaQSykP/GZeR4x0h3wknX/BalXbtnR5gmBDJlmaUhS4PASjP071+yrWGdeePVfZLI9/tyMWl
u2WnCgRhiQ8QcYA1Frg4BBblVjlfW9LJuYRinwUnHFCd+SPzhLCItvJ+06nKuWNqIxbw2v+l/88P
hoABVIQmkX6SIdcEizei6F2bp8UqoL4meh73eO2EOjHOVmTYgf+gD6C5z5I7+Q3mmVoR5mk5QfSp
0LedrkLXnWbgw4bSgUaolx82WcvNV7ULtKvzOxzm5de9qPKoHakV+3tPKDHau5og9X4oaIzu/PIt
D9tga63EyZ69DI5SvRDSBm0VuN9EeB9nwJAnSeYyc7QOn7+u9C219Qgfu+mN8R163bjP1Em55QOV
rd3IlnNJZYWZQg+wTNQcbcNgwLMlxWPqXNgvGdfoDh4pZLiaTAXihJtBGE1fDRmFdgWMj3ZVohuc
v4M421iGvcXTjBkZ6CSsLlehpMuwFgveZANciD8Y90gZcovuxgqC4GijJdOTa84sQgKT6GDUaKl0
CIAEsEaUxKVUggOOyDFl4n4YymBZeh7CuQR9wzh5ctlw94mUGO3H1FONXz/UTFB7BZBHCycIG3RO
sgpWm4F40txCrwPJOLp0edZos8pxt7DHUuzWLI8xmZ8i3Jt+U2KvCukoum/AkIuYlSqUhRxOtCTM
UgnW5lNV/ET1fPBFbv39Tg+/hqvRoV2vOuqZ573GNdZQ7MwEWCleHHZlyFXgJ4c2JyJnqfjR/3qT
YiqBLZNB6sncwYGBRj8HK04Hwk3vkigUh0QEk7+99qlhiHtzW152gg/v/2crONluyzEqeD/F9DFw
Sj9rRNgHtI/D4+2f3fLVxtlvybqSh1InHMecpsDJnLVMKEcg6oZfYBbswXp75ST5MjMeImsEWPpa
O/vfyg1LWwkhxaK9Lbc/QR6EmKAUZuGyyYkUqQeEmi0n/xDpzgL3nSuUF2Or7+72ySD766lwyyRh
YB4+xsej0+HVU1FCGjBwSpvwCzF3Qyh8bjUpE/akor0TB10vNJxR8fB905dfP6Mx1rcbQd/xBl2g
KVaEh1AT6FU3JsHYnkZBsOwYpD0MRy4Kz4dfaKn7T4cSRyHpxgq5j/4F8xqJV/ELEgyP4kf4z1u+
iPAmP2lS1bzMncu2p5fSEkQhKBRtxy2QFpSvn8ZiMHi3E4/IJbPm7oerXQB6liiKv01TfsH/6bLS
y0zVEJqhXM6iENv98oVoKUAJnL3ms/4T/vnrfvDYJHCxisPGZLZv556A0E4tusDngESoAeDKv3Nk
CkPIuh35czIRuLgft4nknUbyIQbl1Gk0hl6+PfLZcLmFVvwimnb2u/S5o0xR4GBrZpj7kwYDFIDh
o3FnirJJT0dbQ+qKl4RoW5u6lA6OkrZMkxuj58j69ixFxdfrZCbOs9N4lj9oNGZAPiOp910DkQyf
8FRnQ3reDYqWGJTE0c/Nj+g5pkfBrFipYmU99y2oR+V8+rlMbbl3po5X+QgTZgK2Vr++3hwF1t3e
AJtnuSOGgp6JVIT9SH86pVnCZEz0fNPIccbvoC7E3LCcSsQlq8FHDtN93U+1b2Cp0/XhjCevz/m+
y9SfLYhttqPjFd2E5SXf4X4BKc1hayrbAmFVDaSmTHIBUuurodcGL3rSnycxHC1R3DCAZYvVkEDU
roKAr97d1bmjaKq54XSPzATESMb8K5jZ9zgCaZbneC/zWpSZ1Kmg15fBVqCUnPWNDiMUAecXDZa1
OL/nEDqwm7BJ3f5NqgMe2zqwxzUvfRILh8EMag13xbtqG/nT51RttRYGC/0UYT1lWczGHDHjigbZ
4wiIl9HCAAcExOhaDduGBE2zBgP94mIxGJgapUCCVJMIxkJajJZemvyy3HOb7d7aAIYB6Zh3bw9f
oLxV+Jy2XJwCJcg/W1f0wddlrk9v0U7zachqTdNzBYXY0hgITkfFhiWIa3ZQjP5F9xDYKx/j8Ir9
+IpRqVKOzJEtWHv5Y4vuZjunGVCS+uAFYdSLP5kgRObD8IDASBtwAkLPYGOR/bpXwaFh7FBis1B9
WaXUXvsPDmvFQYzXpvbF1mFFkMx9ptWWNuNcY6HxuUVFP/Q0bTU4mjL1715w5AY64Gk9RhvHisOn
bHdYuSx87clbQ5wpwWCpVGP+2cA63bysGQeU6yaZtF11vqxcIDk+dM8lGCd38A8l2OXaNyewP7au
EArvfypWPsrXj3ADTFn++YY4+TA5j5Bs6pIRBWCqQj5BhghgewDzXPuB7pJd9catAyJ+wg7EtA0Z
7ySyEZ/JQyFeklhF4xW3FCGWcPJI9d1MJnIV//mFzUQFzmDDTIsJpcI/2bYOGyAmwIyI4GwDfjYQ
xLE+hT5I6m8YZTBAOWNc1aas9s8YAR8a2dJB4DAuH08cP2K24amLQ/6ui193r5epGu1LHmnMQQvC
J9vEViuzdI21RBIyavUNOYrA8DU8KPa0k9/AZ9K8/mJNR1zCzvDG3Wv9NuppDw7swPGl5XeSWF6l
WbBrUzvTEVrWvy/s4Dh2YnZGiKNRjHc+7cP5YBQq5NdvyVSsFAEApTOXmlIs9bxfokfHaKcBr83F
i7B/5FhDPIeI2h0Q+hv1VPI5lxVvE72AHdfRg365hX1hP3oelwggO6gRXdy4s92tmzKNBouW4Pct
fARcV48lYEqW+sZr5hJcZjJV/yJLuSvp2FhFUEUMrS87/lk/KF6E5zVn9ppT/J69SBnVsku9pJ6g
Nu5AQ4mPjcYqt3vs8H3DbEUrJiyzzmgl/8qCjicKL86LWGtaRutoescOtsDq6EgvHnyAmGE/8kzz
P1QKO/nQMC/GNO3t6w52JIpuO78vE2kf5hFJkmjps511xNEqlz0e6b5KWP7nkpaJCZAKXjIqK2X3
1MEttpQ/EFn6ca0wQRF92FoKeISeXuyyFv9f7/K1DNGxByGDpLUU
`protect end_protected
