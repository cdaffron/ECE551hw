`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
a52M0Gdksd4JHYLU9VFmSFELjo43M037tjR2Wm0OFpSPJPc8L/o8DNP64sIaVVHJwODEMjQw0nk7
TRydgBAq8g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iO+OpuhOyeLwlA8MzyBqC5cYmRlwE/F0BC1c8U3pwA+Wv0Osy4JffBEukuL8QwyRK33+M6XA6Lkp
EcFkzCHjF64WjL9ebra1XH2tOEroMC9u12EPPMJTC6LoXhGP28jx1v8BBvDXKD2g+I3TntJzuQlR
dqK2Vizk8Hwewndu5SU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OXUwRneDA6p/uNCdyXjSxzC77GyJFZSAPv1o3hNY4cjOlJWGbzb+ns3yuhPUrFQrpES4Eg9sTKo+
AeO54D7IL7xmMItcsRw+qAtbS/e+CDQ0ogIIkWwMFC2XB4NyVtqytTO9pVrNa/tDhtnMKrxP0ZIp
uBD4nkBZuU6UVE/EQfWZZui+oNHUpFSVn2XtQwv9ciJnbq1Mp72O9QqCKv9eZF32LDQXpwSt5q7n
h8Q97+R75COhvyMOyUihdhOVFIkwj+HdWgj1z0R3FBekA0CtUwHFkqDic5xqh/6yiN+joZZLzeHE
ZKY/Av341M1d58952cq9x5sa3+C4UvvdlXijnw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
No4Z4P5ycD8pGxRsfzrwn3v12+nH419cUxzFzjBqbLSUragWzXgqybjFigwagJ2bSG4+0kd/sjyb
wHIBY+76dD734fb4XW9hmjfhvPQ4X93dpggEXoshpS50PmmVRLIw5DfvYqXQJ4cxukfXfiMjkT21
GHJ64ufQn+hmGQQOecI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G3prrRFfFeBFvnY9Fae0j1fMMJZFUBOWqWR9Xb59TaB5Y+PEXjmcAFFxxgOs0SOIoe2VO9NGxdvL
yS9Nkksj9a8mtaA1y6LRThOvLPNZeWowpunvLbNMmlPo331/9cd8sqGyR2f+64kSEZ+ZsMo0liZo
DzpiX0HCahxUJi9OXEa3Lx9WZKm68G7nJwiDiaw+Be+0EHwOWKNcW70DBAzL6JaW48SmiWbN1yt2
GbKAStox1fB3nqWpZ6XdPSxa2WXwV7j3Pefzj6mSWarGLvitagnxSDnFzO+9wwvQvOlAb9dnQm0V
1T1SptkeeHYKWD8A55cNprhcGRa5g7U4WIEq0w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40496)
`protect data_block
UwGAg4IexXNp04i0pS1KD+eAlKAfxsBev8xSo4rFIZMok99qMPZIAAWU7vNEtEtmK/CwAEsKKaF+
AuFVvG0RILY/+NWFJwwqFWCXqQNGCL0GIgi9mObh09g0ymyg+N/yq569OLc/9qsiUMOWjPO/O3yA
TfgkusVE3C5yUiqMr6mJWpxCPJuTx+7Lt6ZDLDtm4WX3IygSKymNpy68oeEtyZBrMAvt3YcXNMp4
MOTF/GC3+GgQlHS4JLLkA2Vl8fwdRd7ADjgXNozFqo4MdbssZGLBruWfvdYMOjXr/Dfhb4/YgOiP
7Bvsh4vtLLLPFGqNAwRlRboKA8zRsoFMTYpnbvBX7OvUB+1C81aMiWbr8SRjPhBzo+e6ej1rn0VN
hn5FTFbpXfKkigztloqD83lSMWmpUtDUJMonDfbnANXWWfzaHXbS43uS2guDz51Qlo+EVDDgSihY
5p0oiv6WaBsc/m4UudmvCiooeP/DKvMeuomP+vUeQJpgfZagR/LEyIvclgyZr/Q4nbnG48tErMfu
qXB8BpDx3/Hnk8yXodCggvVW/N507+SPNGfDtC//z698SlBKbKyTgEoNbh7ZC4W/cUpGn+ybwTDJ
kGthE8LbKrTlud5YatEdv4p9bEfhO4lEJQwWZGEiBdbkKtnnSg0UlEl8sjpgxSjF9A4VFLpAvFan
GXGIbZlMz0ZwDgQ50RvD/nd0X1g1+ilWpep1F/mm+kLAJzSpLN3mVRhYQMNfOKm0ISghAs35JaNa
tVlQODky2R2gcIIxfkhxB1JqD55ViLTLG2FIb+qbciW7QSZPaBACZfNjdEhr9yEWSKwjdG6EdXE2
rbKCGpJnAicmVfc9zdxzNEEhXFfkLBG39TBzWgFlMdD5NJoim2bWm164Wpf3r6+/SCR0kdheZzMX
rQOZo8RNM7i4MllOHECwUyaq0CLTQmKmjgvPc/Jo0SMFM8oYc6Pev0N7VLKVyxmNf/pG0bff4W44
AmTbazbCLWIVVMCil7K69xKsvj2kDZI0R25O4IWrkjltQhqkN+/ZwLrgDVoLM7XKsD0SupJVr/6x
aX1xo/gOmJuiyvxa2AxXKghTZnad/MitGvGU5YJ8pdUZ87eYly1HIiFQqzB6SVz+cyL8c0jE9UC6
LBRgCb8p6jO8EGVTZtzILMA6VuPnqwt9uQUeUq1z8gOHn3G0vZ0i+Dp/dlCSSzvHUwT72L0yCf25
KLPogevFRuqOQXfULQOx+umiFjdEawAEEH81aYBQinVM+ZSwUC8gA2wIVj5kYbTGZeU+lo5Ck3uY
IJwyUpsqjSomxBPIAWOcSmUXjIkI8vhuyVTTbx3puVdwbUX44dKXIVPokKDrfhBQSb3kksVxMQA6
5hddJz0P/bWuu2Cu0zQPJWOz6v1PSY84qvGqgtmvXWG6LytD1ebmKd0dNiAKLs//xZ6IdrW1ZPtg
t6S5topvYvoqw3MSCBb0UkHxEJ8Dp8vaS9C+Ao3TC+RhwsHlGCxYy9sOQLUyRRlfJmWfG5WK4ImA
EdUUvj0iWiwYXnQpWA9skpq/lm3vFFcMF6IeE9lKszHbbGaDW+z25aNpYLOMPJ+1N6GATcopRlHl
jxE9FZwObaeykAYBEDNLuTLg9YFKSZRNuVaIn9+H2rDGix2C+iFbyxbKXTNeIH1ctfp8ZzC8X8n9
Uh8pfcoHsViKi4p8rSR1IbMRVFkskORZvXyKNpsFBuj9cnGyq6rROEBTwtE8Ze8jGE5NGJyG+g2X
zYgDU5n02xcCTB8iEkikVphzKp3nySgAIw+hmjJrX9nvaBmDnM12xJcumxfHP3sljK4I+dmKs/5z
LCnX3gbg6MlkCgHPYoqy6OdnPp1+YFVlxZnB31WzhfQSedbrZ7rmrrmmC3i94nsI+HcA7qY1fF8u
wEjrLaKFIp0r7zeYcau0jabo+UUFfCVJsYIlr8mvrcG5mORM8NfGUJBZ10Ha5hAjokzQ0Y/mMzTN
0Su0ElUSNLCsmQtbE2iykMixBOX8l/fW46raR7XfBPZrPUfluPYY+Hh1qXVNeaHejX6INJfd23H9
XHfR6wITMFPmrlZCTWX/8O+4YJp/BCcbwkflFdxZTtqssUerm6q67AxsqlF3kwzl4Z+9gVYY+OWv
uSlIc2qktWUvz5kBT7X+tv4d0SzFqFx6Sjhyi5wnjiQlnX8Fh6K2tb8bPHWXrLIBZATRKbCzHcXi
YPFpB3EiIha/PeR/91KVJ77LbUV0743hsEVRrRvJank8AnXj09MDWn+qO6ZoMAArbj0FTGRwiFut
F2Fjx9ry0D0aBRhMKio6Im+rjzVKNnxwXSxAK3ekqzSWpTHo6PJqGLuSBMl3VTfFgALU0tbDqaxQ
6/8Jiw3WAex5vDYsK+f+/qbTI4Q1A77rYLpW49Lv/quFNtSV8K3H/tyB/IxKRjzmfOxnjtS6LYtX
D6gjtkRLQo8lUf3CqvMOyu16qmErzrbO9WutlXwhegN67OUfZ1AgyuADRCp5xCRNzt02PoZILyCw
C7mY6w3pGh8wCnqYYjV0aLt43ekXRHNJrT+99uLQV4dv8FnrMgo31N/3dgetaHjDzk3k1eF4eIVo
dNlAuyS+egJ7HZEUqbwHVVlsvLjUGtJ9xa7IfmmqnAZy0YejvUrZqT7FlE95w41FxOcjcWN1IdQh
Vn+9AOltx91b1ViAudEkAPUrt9W08GIhVXa5JYD6B2ACZbEZ1cqViQNQ5ZufXBWa8VffFQisKjQC
qhOWLUTsFPbpPQC3W3RuaJoanhE7cQX91M8ePI7Qfd2Fj8Kl3nNup0ix1X/C993j0SdotrV9OTJq
ohrMw/aG8DOjIb+SmWuaYWujiASUv92aqmchneA+Q4ZzR8YSJ7aUowpfNhx2bdIp9j+Z18w7njKY
XJ/Kj6D04poiQv4afq8LMlITgtobO5wfBtJ7Te5zVE7DqvYZHE8JP73R+EOBFRHtT01OoFlT3BOf
wNLk1JJpIZcaiSycp8HyRA8Vn5YdhEqSmIt5M6gv9tF69XP0aAwk3iNV8UNYFxxfWn07u5KFniiD
8tms6ZD2rCL3H0CptwHtH1gI4LJUxL9WUSrUX4s3p8H+QikjyfOivoMRtKdbNAdCzHXZ932DQVQ8
L3o0+JNJwEPyq3O4PxjjPokvZXZkwTHPpHvwhbmpJhkFVAvDfc7xGy75ZqT4yahNxhEJsCxJFGk/
lSHxFx5UPrCFJ13KjTVzIX9nVMjLIldAvTP+jkHKUeqEQ57i3iJJZtJiXPI6Uwds+xvUL3QIyaQC
VLM/W13ZGQSXBte4IRQkT4e6TSYtYRc4fVtuAHzfodhqiSq/QUgEa8kD460byy497t58bKG1VgG1
YULRujxiVhAxe7h9AAR6gA1BKD5TcEBVXLOXJHPH+Ufe4V6p2yocMeyW175f1Ns3XGQDO5bbv9w+
CBF7mIQegEAVkLcq0y9uJFpeSa2bQ+mD0dwFYz1effi0l2dFWvxmFYcEwArvodlQLp6R33z81Gkp
BduIR7E5m/rNUpeXRUnhxva8Ebi8ZTp1wZttQKHlJZD7G3F+ShbKI3FgQ18gt4aBRB+Td51IUNCL
YP0zIlGQWUhEJfNXLGotgF+ht4jLobc+MyKgjRP62AKnsRypSY8aZzAoRyAdVMmluJJyp4P4edi6
BIcv4CKnrPmFrIYSt+davqem6hV96nwFEyzYa3FBLswmcAh8LV2ml2MW3/Z8ozcMliVVgz9swp9u
DR3yTkMTNakFhJGt/e/RL8rfjENVxzA0nHNdFuLpSkAeAeZ+dyE/bVxB4wU/Vg9TdVxmITilZUR/
afijn9Upxt0NOMmTHWlKw58LMgRCk519iyV5k14qwZQdbUSNHJxDJMGYKG4gEtcpht639agKD3wW
xZRRaNLM3pVaUsl5AiV1ER0y2e1fKqn5UwF7nMsJSk8tGiO/5TZhrbJ8mMFnxX75Ay6SOVLfV0ao
e/xp/JJjpo+6cKXmfx5aCj9bPfRWYX7oLkoA3Ynn988HHE0SrU8WzeVoWJGUerysp1QB+CrqMU9h
/shHdLCOjDL9kUPjyI6Y0hF4p5BfHvr/vk7f2LLVJ9yieU9pWUtPmE489t0hEQxUC8d23G2Hpqkr
duz6aFL0d4kFBhFGt6nSUFkJH9jsdXuzVcx7PnHmNefbbdZYngkDN+1dIbo+jFS4p8YJF/ZqYPy3
umqECNR9a82Sr1DOkACA70oVwMOimh6AEcR1vQnHWKTq/uoA1sO4Ztq+TLha1Irrr3854n+IP+6/
TszxU0cFSuadprQCqyoxYN1eOpgv6vasZcd6vJMGjeKNrS1NCSjp+KIF1U1itgBAQLAoe6MGccA+
ah+Qh7MnX0s5HXz0JpodH1ANmjZIeL2/zbbhMUuo8MOgf4AJUITYuFr6tY9boeYHGyb6UNhjQ+X2
L93apTBQ35I4u3/IRyyDwSgqVyap7pNZe/JNXXiUnso4iQDYEs5SsNyNBMes52tbjhw3aNkp3qhN
LguTrXPM2HgsrkXjcegKtpi/iN7b5eF5iEbfp5ZumU+GHOoNMpZZN0qZOpTeAePNzRFz9feaSgMV
KUgBHZRgiiPd+6b4Un2xQi/YQKiUupD/iDg4VlhhL5+C0IHjfYdmZ35EJpvVe9S0XFlOSVNPli72
3O/xavzCKET8u/PdK9FSuPdn5A5aql8Gqz7KOC1GrtzCJkoxlyEHNkN+L4tPavIHp5D56PBSNoYo
qd6tmFdo975jh4147aplw32svHEtY4tBW7FONo9AV61bdmbDkElwK5AUg7JTMKTHQcswQ6F7UYBE
LEGza6URQ5wKFgkwndnqGdbzvXO3P5CEcxwJDURm3vfWGYs2a5mzg5Z4yKk1fWVkO/+WQDm4oO1b
C99eRMDRJ4guMpmN3FcDqpbAIkzf7gS0Ov/CpjH6E7r2j7p2T/vceQC+WFrz6P/oTYnjBy8L0rri
+UyT81ge2e+B5WluzGvckm/HaV3OEx6r4lcvm12djF6TOyR1fLoIEmLki1CjYm8fqiOYAzOPuaMO
dbZfPgFD0n/7T1JFJTBUVthzAoOKegpgK9oV51s1I9q750afDo/6Db6nWg17O4TjBv8meAtwf3ye
9xgIWPBpR5IZcR6gY9USQg1xtZ1nRIzU5nACaD5dx9ScDpg73aUVlIFMAl4INE9yisvqAvLzq/77
tuJ27TesxO2m29bM1AWnI0d+zX4/L8OyXnqtNxylbnkmRGZ70U+sz5SOzWVWJxl+/b0vkFbUcFX1
0TFqDEl33Ur3v+PRnQ2gx+4xRgtewQZuEw8X5xkdMtWjGxqLvdIv9hn1z1L0hXhihfZuFGxeIi/H
O3/UFn07nKpIrfAeFR0AxTds1VRzTFH7R4oISeoKj+rF/5+GrA3nkn2l12+yXhwWPmBho49fPKol
64vqXbKa8vvlA2j8VoymFe22Pibwc4x8gEQVWQbMCTGU3NlT2F5mkz2PynQmjnR+8n00PimhKEoc
Pb/u7l8ABSRaU5F3cnH7+pcykZ/takPT0NNTIInBDc/vBMiqFR5G6Xgb1ZLHduWov1/1GyKKI/Yo
tT3LZuSm1TJPIRLd363Iuf86bXMY2swYrpJaY47pUAPG/P5FBdt9l6p+emoxQRZP0zvCX4+AuKqe
6Qaq15Q0fUmrfULBgzM4DMQgJ8f2E/Z0SRQFxcyfjr7uiN8dIsWw9tzfabJZc17gHp5J1UjBYet7
XsYdNNBnKnIgeV7Zw4OfA0ICmeJ5nechzSJwpZU+jK4dBgq4StVM4tFjaARzotfJus+25A6zyST8
qXvXAGQHY7NH+BadzX1UlNtPqPYaoDtsOICDioC2lgFSzC2MNfpQoiWkm22rYKPRoEhUmC63MsFZ
Z+BclKIxFFuFEZ8mnc1MYOTtjfRPF8DYsrLlNk2yh0j3bOuMVWoBllxAvX5dqTNVVzf+ArUtA9dR
oTNcTlN3qZ3ERcEaU83Qmv6VSd2z8edxkToOKCMaEkZs3wWtb+fysKKYSkxEoNqPDJJk3hoiJ/L+
Fu0sPTI1Tshfi95GBghU3aeI6//LtkWJw+Gq8Uf2pMih3XF6wap15d4R35IrQ2iypqortkG4jgXL
IgmJE0/EaU/F2WAhrH9GKjwMnzmzlHzvZLGZjobuDs1uEs7El84hyrWFbod/ZPy1Gn03KZRmbU0E
66upqaHg/PSQXyMd9fySO72aN4ghuc3c/1FKgmCsyg1OxSppjv3+2Pigw/8Pp5EbBRCTO/BfLbZL
TcwuQCoJJ19QBFDUsoRb46q077egVgNc8nlLw4OhSOnqrX2hvx31koYpgm4ep8Cn3PhacAs7b+Q5
tDUjpLFlyNIw/jHm7ZS9nQaYTwCp3m5Fp2lZ5xTBUThU9aHdjYeiBAUoVCKQe+aVb7nbxlirTMlC
OpVKNApwFabgMuFIWKb5+s9w7k5UsR1siVaEPjak9Ty7eAcsPaNoQmSNYxpC0PQIql1q8UYj8fI5
Q48ARXvBpm3CHckILDdbWuIpu+qjuD6E/O5bhxjNVMGiTLTdwlhezqCrSYZ2vACDNZztj2xkQtU+
2logCPVm2LhY0FmbKh8wNZEmB/G8kUh71dUISSZEohUlh+9gW+7FPRnnswO1fJUKVqExrJQa57+d
wa+jvXhRmIY99owdSFkaa/Uk0vyj4j06s3SHxki8Paz/wy4/XajCGpuPbVsTGwunF7qNqpZuFVU9
FfDI9/JFQhTIsNhytCBffhM7L0RZX6asHPEAaGZ1Jpy4Q0PWDDDXTq818mU6wvk3vgkmUdvwDsLw
YYJzuyTJ0Wd5SlJ1owMDs9UssSAC0b7ikIc7zTo6R3VvMAOEXIFxKpCqYj06lp8pSPnZKcClD6ZB
t6AClpRAbH2lCcVTCh+NMwDj8HAw6ByBqwJHy+q2hp0cbTT9B5/Nwc+8Xz2ERJj20eGPPy4Pk7P5
hT+6ao5wiIhz4y9h2SKFUUFeILmBZxl7v3D6DY6MzHCgEQxybEkqu6kNdOmTIQ1DkvdB62nyofI9
aTOg+XD87EN1B5qmU8FpnJPtOrSni/uid/DX/HwAAuuFXrj1OWm34JAvNE+BMnV88fnNe4NKlgBc
J1zQbdGmY8WAVxpp+BH8gC4jkqj+txuuwiei7sbXdns51Qjk9HJoB4JnhGk0psXk0pP0cTJvhFkQ
yX7cwJw0zXhkVySOBqFqVf7OTql143PffLflewzZK0R+FM0Ecr71JmUssv4R5tF2Pa+attWTJnp3
+bNLniwr74hLhOYKpztMWHbi/watDwY/eEY2THHwB/27tlC+HKB2/sWbEgcvH6RIomlZhUoDGF9c
gS+xMDJC1FeI8h2ujDolVm58zhiJVavKaLz4t1LvrZJhvzXo2vXKsqkZDNAxonbxYu8r3wwTAwqN
z7ghYzYl6AiIlnxtt1B3KWBnBGu1CLMKstGbZ/gr7Vpi1Dtm8f6RyTWbxhEgwT4eaBnJS7mXXzac
Yfy3QgGHsXgM67DuhSEtiIxlAMWmMJO5Vk76a3bkgURVBJDMPi5tBQoIstK2VIIVcSWmC64IMZai
4d6PuhtQ1JjYWsu79ZorSING7wTu9yawIYGNSdOEx1W6Q0GycpE4wADzXSludcML0NRX/KsWLN4y
vQXqeu3qTyzhkzyyUJeZ8pSJv6mdZQ6A1qJSaF+T5iMWLwwmnQNR1m/SvMKFSsn4NF2LSB1mWRwV
OL0F8MpRB4Z2BVGmQv80PyKgIjU8xuqr4KcNxJp/oBeKTJdeR9Ro29l469Dml+kbkfDBDJpb4boR
gwFlpFQGinI7KlhqNJZwuWB61oL8c4Moh/o2IBIwWTO6/4NPznjxplE+P7Auzcron4bfq/2Y9tZP
YO5GkClUG5AUU0sZanyRsDXLpONbMIMFFvW8fGoRqwrsFjj9R96plL5RSeE0WyVXCYnOdr5/nHY9
drD6BG7q5H7yY3kh+Q2fEQIkfEBgoeUVaeyyLInJGdOwkZWbivl265tQW8dP1WMzNGp3tOThZFdP
AJufziFUuyZh5ME+4HgRPoLbdJeRMBDX0gjLg2Fm7JHkm8Fd5K6SuuHKoKOMpfs5qbz96hC3sI91
ZSOsJUMEF4NrrSMwWjW3u3oOqX27UbAQ97Sr8aSw5j3HgHe1md1GX6WDjZQEn6shYeEioqSAyMQA
eleIJr+zXaMJX7+sCoR30Ee7DcBd3TJGVc+gx97pz2/Lr1MgRP2VlKpUhkA8uEEZqOQsrGfwO2uw
trSfbIiiKZZ0TGENbgqxysYMHa++9HQtyVIVsXWJsDk9s/kxjnw1culDqANU62NfTJ4eN9KsAvLL
terCxH60k9gIcixaCgiqQBR7zwItdMiliE/iSoWPG3ySlthSs6LS93EheaabBpeaeuPScuNe5UCM
ch7rPCKCudS7zzEjvLdMj5122g09sBsmdzM5KsGgvjXWGw8pyymwBZY3NuCQ11Qq6cHb6UfJp/zF
sGp6b+wCc0tm0SLX0/N3U3lCo2Z7WhLaOZjWhZXE3xVopkofRa7clvvcfDtQuazBhHS//+4j0WWu
SNMVMfo4KKdbCG3sAjvDRSNMWnFAHRwpJRrP5ti9LN4gOOuWlSWcvXRSoyVR1np/W9YR363MN6Ei
snkkTzcY+JWR/AcTCx78RH7MPwYJYBhW1rHx2KtGX9EGVZYeboEr1tL4mKIlcWSI+fJh65MbwAhD
uz8Kt30L/hBgRjTYjUoNc8ccRcqJV/srdxHhjOf5EYekHbPl0SBVxQQaC2u7eAEXfEAg3LlXuP8f
cCTXJkrbqLP6DcPpWAa6RJIyUCo39UE2aodbmiAiGdkjtc4HdVKIh815AOZzaOluzAZiuALqrkon
FZKM8Aexks57KyGl/zC2ah7JiLWyVTE3PsTry/ejHqHZYIIHBJUCIo5vRXGUoS+umsCtAuw4auWk
3efg+dLcPV0oDfjf8dh5dmy3XpYgxO2fVm+/xuy54j9EVC6voJiz6d3TSzojhf0dcEFisyE+OBEM
Ij2sYjSFdknm3/IQ6TbPenbFyvJanRicC5pEGt35Nx649DKJrASOjw80UrzwxIpc7dgwyEiCHGLH
ukWI1vASmJHpJF0SP/RoxkUX+7cUc4Ap0OuWBqucU1CtIbr1jBjlCJTgkILoXPrz/NKrich4mM+L
o10vIox0aiHD3CeGjTz2Fi3FPzUJjJWPnwB+Vrgfu4oEztRtOEj2jM0kQ0/7JKz/QVD7ixZ7nLh+
Jz05JLcZo2etFikRa+Qy6CGbHPFHJX4g+UJT5KI31d3EGDwo/H0J6lax9QVxjrvZipG6mkUrZPSS
HjrcfAE3rt6lcyn3/vIZpbwlLl9bDAI3SYhDPwEmgALvmxspHIKM6Tcpjd3Q/tyYq78gamO9WhgB
dP07sBh/LI6sUW4Yvj3A19Q/sDrFHoxU1pZjv0/r/YwIxIYuDwqpKsuUyVdcwFNW5ulge7wIp0FY
7HmQ55VIKEFRK4YGdBOaNKVOmj2yfc+9GpCudOPJWPUwCBoRR/2sM8Ui+y8YElUKI8pPBCNusP08
Pbs6DMaJJuB/jSgyJ0GemTKqv2jkOZH2JKBffRD6Ek5sOY4COuR6a7Q5sAo01rX+548gHPigTvTV
pxwm4nPcROssDiUpSfnD9VfVl/FwfwhMwWZeSigNEPkVdx+BBMQZ0aid3s2NeHN/gA+boJADNcVL
cwStrT3jtpzPynj51FlK3NVK2hHf2bCrlBsKWhxY8aZPlUoYXmtptgfJ3tdTpqw+8QDCv1cdIyO4
E1GWJLnxqzikzXpQcgjauRwWtVpT1S+Okqq97oVGh/JxyTGWsgGmtdmSQtCKo+gNdt75IhdQ3kl4
0BAexeelwreiIlbK+xS7LxzNTYZpa9f0PmnR2gEhiFBE5ooC8CIwT3wnQnFCeih7zXvpYFb1NpR4
7BjBe4Yx43Q29eVT6l+bNzTxe3jUg9YUjVXYb3/a5HVN5TEWHAIYhBfi3+CPhg3ZUTCvAgGrqeTr
nQuE74Ko/wjKRURyB9N5BbmXx//ehhigZrIUkClPeQlWY/SRTb7vyKKge3g03AuofsuYu7U45Z1x
vhqjH2Gw9/1qz/hw6VGRRvu6DrdlJ7N+VvOPpWZK56h0nPnKXN27ol23ao8h4fWjIZ2r5Ej6ybh8
vpkhtwsmUgZbh6DlxhPrbmPFYofZZsr2QBQcRH5NuxBZYMLOaJIuASM9s9O3pT50EmKH+wns0HTf
x6sXmjCNmghmacpI3VJ7uJGjF1ooDTPNPMVhmPyOE54jrnZB4cOV782l8/UKyXU2W3hMON/e+1Au
MSmfdlOZCZ0M9H3qZoTtR87s80SEj/t4XViaByx2sp6TGUG8VXYzUccWiC7zp9RNsCXcdmPwKrAX
Bx0AmYSnXWu5NlnrA9DOvqQORAQsg7BO3/ZMPjI8eN+gY8A0hz7Qz/u/v4H2i2oM/BZpCCWgI0fO
VoVSt85og+KE8JHQhy1/31D6a+kfODLtxkjTlsXYALvyHiVT47um3ltkJUzwjVwGRSDwSzWplELT
NssA30WdM1wSwtS6ciGVY1IdZ9rcEqkUHZYowBj/QZblIYiHvmwbz1ft3defrRnGirnZ5CM0bq40
hC8LrMjXll3RFOk5dt6NwN225QkpD1pD/m3KUT6bR7ZvNKD/L2RZ6hyvK9qu0/0r7zxUe+Md8y5L
huzGhSU3XliAIMkXtLPG/28x97lqtEVlMKM/dbApqgWHRzEQ8nO6U62mhW0mtFt86Y7s63dHkLPh
mFBLIoatvo1zczFjf/uWezWkr8DFMfaprR7zX1GVuCiNtJtjrkgra7Wg+TZonMoMp8aW0kcEf8Yd
LixjbpcqFOnRji52eqyQXtcVUtycGmj/mar4UfOdIazc3KRe2tkHkqoNha9D72dU7JMOirEMwL9F
9riMdlC8TxpWMJy1tW69980ZFc+ZxivK3BwVxTAE5d0HPZXRdt70exDs0L2vWHvG80tusV3ODZ7F
o6G/eKIE9G8/E9E7oJEwtIAOcI7uqvb56Fm3aTmZ7cyEA5WyfXqPMmrAPuZgFqcNK1AAUrfiq4sV
att0sOw0NbmnswNv7QZkSjKtrdhqj4jFZqq0E6+zWMEvdihIqsko9V4JX53YkXKtZ8zWQbVXuQao
+Gn3EKgE1qpxlMJY0uxZIsyfCcse1hBchnVslm3fTRiv4sOx1pEMerK5yoEiF6HGOK1Ag/m4wAU6
70Bkv2iJrhHxtk725s6CBO7yjTFmyWFXlg2jqAvtWr4n9GbjAGLdGE+xqRAadNCEQWxvBW+4sIgR
tNGpwpwQbCswfLbjXfU4ZSPjYCO5cGfUMfZR8pWn6JZ0kHqMo1ieJtl11vyzvaG2bZl6agWrMb7j
JTh6wPlu3PVpzzt/nCkuaOBCQLFoEiVBOkPJBaUA3m71DjEk+44WUaTOirQ65UnUo5Utp1uwjEKC
eXAg0oKOWJR70JeSlkm/CIySMwnQJIB+ZgcjQbsnHQrsLCRHhHURX0jZZ76KtUUkJh6KHUfpOf71
g8kM4XE853pR4fhITv6ulPUIR8Hj3kDjUXlpXL4lgWqpCy1R6feCL6YtvGrjfSXWfT1vpK/frYs3
CAKcHr7Lc04nnvgSPjxVN9ivuyzKCu9henqbB7yHv7dw5P4UBXsyIHT5Pcdo5YxReSNSlOC8bmAB
6R5w/7InOc/6lHAa3TU1gFWLIg0h3WNZAWH+hC67TVYlf8ur8afZcRwgIZaIR0wJsVB5vjy8eucU
Mh+eU2wcvjx1vjIOD8ZGMgE+EGoPZlhOB/v3hy9S0xDG4uE88uOxRJG1RG3/q5ab6jwdn0fO08Jd
emlwvRreOmzWX9upeIqLoSXk0kRISTFZy/UQysC6pgR0nDkWdUlw/NgAV0ebHpXgDsiZWjm8JwuH
g87ljQI12d3bvdeGlWyxa6zOvuH2eq2FyVIoFc5Yk9O40T07KPGprE6THplC8GQdXxgdTRxuSIlC
az0GCBl0D2QwP7/2iJDHuO0AOHtfSYZlPVSM2NvQZXojwUz4uzsrMTCMdSlqJQvGV/IlC2WcbXhX
2N+da/5rG1LpLLjrd0zLiSDgJ82nxwl6ocMjjWNELFbDB6b/EKqGdWWgxzaKhgEM5eqO90HNeFYV
SHWcTJafcWl3midZWH3bF/P28ngGD/VKLHfH6LwapsJRzmhPRi4RIRMnbsYgnCW9DrpP5dNQUuEh
hUqVvk76KbishD6RnpWfKt9YO08g3io84c5FWVgtK+h9r81d1ld+R60IizKMw6yhZYsvysYiweI2
OD1jZBfLI5CbK+0QKds20iHxXtj0ihP2g0wfvj46nP1P0bjiM3iP9bacfIOHVglnXMkuENU8CkNn
MBTdznrN0CNPzGdSe6LHW0c/zv9KeSaH1nQUI0I9dzypEktFmGs/vZlsWa4kMRtt+F83/d7c1DSu
ukSdpeL1mXqgyF5vQJ+D26vBP9vD/M8uYa3/XFF6LR6D/xaAubS+FM/W8e01FApp+S0AEwAKVsXx
9j3VwTSsMIhi1ZjZYKmirReWcrFixSI0K9itz4Km2nk9Cow6PO2zWn130k4vqA6O+f08QngBZz52
aqXBiv4n8Fb1feFo3Bckn17FbY6p7jB14ilTnyfW7+57ZLQGRWkdLRvxnqa5RZj4C24YexkhWM98
LgEdfB/9vzvC8utMJmCOHjS4fkDy6vKcy0MvxYwbIzgnY+A3SuubhOKmlTQdjqgp+dGmKZhBBr5H
ueWZVKoM9VGrc64yeqIAJcB6apCFE+bjXgDOA59dIQZc1sxcDjykHTiVp/s797vBRwQFtq13893z
cuHdC9hLqKtRYx0d2v4dNHcfTsUYHDPyf0LVVMNaLbpbv87OFqyPiXUzmudg7Bq/qhqlIoeAjw2U
c+yhh41/crz7pIi11ZIKb0WpFmUkOSCeouec3ziXmhwM1TiWTgrb1GCgzLNPkbDhom82I9b/jAMK
z4Jq3lNMODt/QA/FxNXEx3sDrOo+aJu2djMXlnn10AtoIoGLP/eqMlTBu8+coa6Ic1WZFvrfzrxn
EnqpCBsClY6cJ4gQkcUEDSP+xSPT7WUtSW1uyRuY0AtujrGKsPERV9ED6hm8ziyDkLiXRDSdHC2v
4Uz+5NN4CydVuG0SndObNZBolIqIdWpauolGLNRrSwzum42LyLmTWoaRgYDemi4bxXAHVxXfvdvP
VlfYpodalF5wliBKu0GmOOtsJphfXrvLqeRfpmWW9TqxYrmF6EmhT26dkXKBfFu7KBkIIwK5RpRV
CPdOT4F5xcN354FEcw56bfpL6ydDy5tgmQ0d2fF5+Fr+D0nGZpK4tDJhB7wOVjsWYS/H3TKtNgYa
eadSax3GMNAidSKQ5HEQWAkoMt47PqC2bDY5LBp7Mgu9+x2m5l+8He474cuUcdoX/81X9qXw06nb
Um3VALzt5ffTi9p2/agxEgAUNSb5ICNrF9XaiDCu9DQ07on2iF3Le8JXyEkaOQ5W2wIHWfcuX/+e
RMhOI5o9hG9acOtAOAxa8rLfWDA/SPjmvA1tPdlW1uevR37MsXVU2jVyEPz5rhv19sW0EKDaAPXX
GLBL2NyDjH7gHld/OoEhYRAKFQlqgIHQ9ANvOK2JgSKpH0U/VYjhD3mP7Qgottv8+Ey/F4t9/q/j
b1mdCQFCcySLs/HDyiRkADbYxtTRg63WeyPSl5NwvvzTxnIGIhfP3CmB4miNIm7Z73mlMz4clNeb
hxd6Kkr34QyGxd9bQ7w2Vbz1h73LxDkjqOo0O/wDgCUsbQeIiBeDjpNDPalXcsKsOvmDe6g6g3pJ
55tyXHU/6ag+BcbzVi8bWWKgy+yXD0fPqQLL8FKK2bqzsk3415J0EUPJd20SUzt0dKS1vNolK7OF
1wVfKvPr5tkl1vyEpFjBcle6Nk9OvGSQb7ftmGdj1VwkXgD8ashLc73qSyMIYdiwh0vPMGnLdHCt
YZWwSkdZKYruqMG4qQi8+K/vSgHAQr9WDtfa1QScK3uraNLwOmv4vVTbBSYP/mz8/zVG6wYGlrYd
fBxTmm51ZP58peIWH0kvsSO8lu/JLe+9MxQAKtLMgiUsOv+OQpW0+IIZI1sT7VrD8YDirhmABgDD
MLR5MsuDEjvGv4FNr5InNyAsdoT+es8ZIpokH8e0QGPtDH5old34cIQUAcQ/Xpt+GYBDgTdnj6D9
BEgsi/egtOdOeDOBbmRpFBVl1vtV1ZsMwvsU1/OpmsjrZ+pMNXluSp/44OzmS+58TD8nahNCIY0r
3OSpVVldoE0o+i16z5U/ILf3Q6qxMHTg5NlT6J2HJmQhwzk8U6sM8SEJOUuRGA9e7nAEclMqdsf8
CsngX8Q3DRqZTEQrm/oC+dWDO/FxZ4pjxBmeeESpRN4C3MTDMgQKhJYGIDY+wsHPHcesYm6Sy0AH
y0L9tCs4Re6M709cHqwEfbIsdItsIhczTCjZsYO6FH2VD2rG3e43HgSsLzclSXsc7epD7AbjHjLK
7zp7lxg5uh3bwXaHyu/sUIpDHpeXGJpg5wGZ4lrznW5ObiMdlhyBnraJEkUSxdhssYsRw0NNl3F0
j1kXA4CtT5LR6CLOGnsRLHol77i0y9KDh8aSJ+RQIjS7Rf0vyv/kQXPL72iGZGnWi0whsHSb3xLs
DMRL0PIacHpLKwrAawB5w9CRJMmOLGVW63ccpoN7h0zEXsKsgDzBuQuud1eVfEHKU92rujNCnfDG
+GOBvx4cdwX9VJx9JxC1jwCGWkgVioB/mqbR4OeqR3QcyCzUWC2qYj1E6Bptamp6oNlak85R3lvZ
4XvANusnP1EgeT9q/xLibPsdRhss2If9dpA9uKt/WLORYlj3mn6SX/a9sWPj9Fb/yO3qX56IWfG7
d1cSLZRqwEy204pY7j7EEU9k0aSLA6HpuxcyHEzEYqxfQqOQt1RJuI5wWSG5SptGj3L8ZhHKZzF2
kb8dOcA6ANHG+WlnkQexOP3yTxCAKO/gykK6YjNBB6ngz+MlpS8EfOY/4MiLRB4W9/OxJr+mD7J/
kFR7ODie0alBU0AxQEjNf+gHR8/G6IEgzofNPb9WtZlEQnczE9GDvC+gkNqX49vC7yRm39/cbwCf
TwtB7WzhL87hCgnmI0ICrTjdHCg3ofsHg9gopQUojvn+L2FdteuhARhINjurX8jEpIQ3EMZUtexC
inTt8cf889C7DzPqF0vVZhnyvuBovVTkInfc9BI4UaL9v1Q+0iCkR0NLNz6ZaHb1dGYfLMkDyA45
aixIwUY2yJSke3DqocJla8DxK+/Hna/oArb3Mh7/L0ZWeid70xIc1qkcwvVvqJVZHAgNvtRS0Whq
JVZLr7duYF8+1q/XDiYOojTP2ZgBpALEy87UCzyllcA7TAWGD8O0qFtpz26tY9QOuoVhhj0zEVQg
u7WShhXLxAhEEIFZKv6TO41nUYpxoIRY12VGM+nIbaQBXd1YNzIFEwGGnsYmrUA+mYGDkNd2YdlJ
ILbRAOkDIfnQQFBTpkUkdSzOiMvSTVVvqWvXGsr9BJojFs0ckOQtjfMx/MyYJyszzF3+EtatwcOu
I154LYsGW51uroBO+KIFQ+SPpeihfcN1M6rMfPXh/c3tvHNog0SIrv2Lbya1d35iCdaEMy8LeO+u
SomcGHNkfWjNAJ8OQU5suJ7UE+TjEmXngwAejeZ16+VPCl1gbAM9pCZnQ5AQh98eBe9Q15/H2pXm
S3tLIf7mqc4uKGhEPxeX8QsXb60a+SGuZ4wVXZlco5gD+lq2Pf1ewPrvFx/v8iYINwUmQGShMUGX
/rdN27+XlMr/kKJ3mrkA/ETN6P0Slg8kLexCUNuKlZan15qGF9bpaHZ7QhchUqEMmguWxSL2HoWJ
OE2d4LUgGikaYgc7BxLcUT/KW11fu2sdJGxAUZRwNrG4IWI5vOqT77/2kOA0QXKb5dREYZo0jSHP
Zuo9vBdRge3MowGjIE1AYbuK3cZjaV/dz5nRCnGr+RDh+msPJ1CTY70OAfPsJCPDlQW17VzkwaaR
Istt3Ux8Gr+mZ4csh1Gd69KilvSbqi9eH+gnkliBRFoM8prUMZ3UVTKvZXq3PeYE2Q8CoZ6Alani
myh89rtWv4r1YK1RIB9biDsRhEWvAPmZuCPeBmJyQNsN7OFXjjKKbF93IJpzoWLYIWg90eqpYb3h
8nvDVlxvJ4UjQcPvVAoJmVS4mhkD/buX6eaWugJIRfP66sFAx3GyZ8iKubbOmH+jvcE592N8fC7V
KfeLZODDs8n0OmpQzSjI7iavC/xIo2JbsgFw9A0gL2UFhKeHlfWSZDPnSZrkpuwCZgEVgtcgrEHC
lQWGqa0HKNRBHogXXUXZj9PzYES3bEr3QiRfHESLWVHCyv/SQhLVuWuI8GglVEVo04Ms5uLCAs3Z
K2yCKNQI9kQl2ftLRqRs7ZSmfuBhLquGckc/bdGCSiXzLKgCKKehB2m7Q2659KlcN2h/p28VQ6yr
mvwe5jCeIyhcKjR1ia/j4JMxiG34oNBSlb+FTdygEDw0qIwlv0bBpkLdzbK8JgMGNAD/pWMxayKV
rk7SgKgLwDEt+0YZskCdTYKXrI/bLFtJfcGv04wyLd4Q3AuDyljZIlx20hTimC0FMh1Y2tnHWOXX
vNXu7FrdLbHpMYxNeI/FzSoqL0ayypEvxa0Iju8NY13JwA895Dgd30kH7B7rEi5OARD5HwM+BrSx
IzOCPdpneXQL7anL6fXukfuoDhmV34JIh1yFpwOYsYYLHGloJPskkUsykWAx5ZDAKZhbZvV0F+Kg
DI41EKIOdmSIJIxCTpI0D9eKhULXyfx8qcdmOwqPS75e1tXidcZLnKeHitYmbYsHBoi1q50FZhuV
B8bDqDpon96VJ08pwYp0ZP3exEuewFeVeBBHEADzKMG2rvu33ftzLkQuqMWPPkX46BR5cR1t2v66
YjPci5+L0QkpbXubmCnUn8TPFAJPCzjYAIKaTceMvp8XgVDi8BcidhDbRNsdzkMipQZXd2VhHtpN
S6nUngAHPTt+Rm7DT+r9lhyQsI8J6Sf2QSsz/RLMBpP+txmJZvJbvoEoq1HDP/w35slGMKJ4NlnF
b18LqC4sv/Od/aX2WuREruu1hTe/qpcw3TaA3BnmZFqgkfqokNq397XCVFPMHEetp9I4s3NWEJMd
0EQkGazTFVlFkoHDqDwGny8sadi6o9clr7niv7h2pLDUnprl2kGi55wEHxIqh/4uO9HrMQ5wtH6v
fpzl508YXX+PXu6PYvPcXGN80eW9e0FkBpqPgF8qk0LCHWtNkPeG6YWPg+rmxMTMQ7G1yBdWvnR5
Bp7TKn4JVQn41v08dcS8enf2pZKd873OjuMtD6hPqpS4v4OXsUhsPtj05Kh0kNIqHmLGQwbFtbYY
zYDh5JLKXKcicWc9AIfRlXUlU7qOMBs9MBpIprsDOK7NKnzVGK0px0DiiRwXx+jhH5WrwQgyPqtV
zQheAysPQ31sCpAX/ok9rZIJE0ThkI43tfouJMjyyUcJxE81Xg/7KBifg+rZxdLPkk2693Kb2lLw
iRhoexczfOephJYL8ruv43FEq1NmBGQj9Do+J4PRlZQ0Z/YcOCidFmQJPeEJlG2e7fwzxKuKRifF
bzj6qt1GKlqRKPKOEnFV89vpJPc7+6jKKWUkyk9BfMwbbBjyKXJExWLM+Jja6wGR8GjYhMbs/SL6
ERl4i08A8UxENwYXldoTYGAJqwo2jdMaiHlo0NU/B4VWW7bNlOOSodojRxxzvu8Z95TCosJVFsXp
4G6RBhgdfGh87wUcvxbzmsEpGnCoxP+o0nGabj3Lh2MSLtQbp++k2P1snLZaOdvf9mWuLj/LPMVd
kQOyRmLih1dHkW2nBGlcQoXCGcGlhOl2mt1dT3QSYMLCu8BhB14o/JCGKCFNscFAqYAH0h0INNJI
IuZxPtXS9yp+wi1jQUlW1UBg699JAO/bZaSXh5etvgIMrnUlzddTKWPM8CTZPeK7ksNOeLfTmah9
tmcKF4xaFlJnCx/nrXNwC2uRHWUlc/CIHU/raPQ151HrzPryWsZz7pahfpCJBvlAM4FRRib7OEqB
HmnJtn0lp45jcdauYbiZz86tXvzIJvNf8X/QgVGG32zfSXXZ0ptF3iZjkS6FFqzQRsS/2MbJNHVc
S3ajrbJ1ZkeQkCDyrUSDE5VgLWuh+249dWo805HakspkT2/hUn1Suc3ebJM6XzsoiAOu9pnIWlJ4
+0PBWnztsYhtSB+LsGaAKLf0HiFuQ6+X4hropyNJlP0Ct0oYOir66GggyTyag0uYEGexIahWKG0u
2V8d+AuuBRqnsl3p2nNnCowuXpWOCkCreQpNESBHjZGKOlLPHDBtrsU31qvMr0F5aVlzgQ2Bi0OY
cXeamtLE3y4EPJex97HSHDqO242kteR33+xqjhsPIwmD7XIFpKKGAPvYKUfHnLMygz1H7xjsax0+
a5esPm2azERlP/63oqSBYzaYwKwIlvTM1pUQEtwJlhTJNCudNQlYCpFCL551D4Y6ZwQmWTo00EQ6
fBpgWdFB7kmNupp72pTPuoXAkiLRw2tbcwOedkbOih1MZiD52x8yUUs50WyovJN46B2fZJG3QfWv
PsZqqDqgPldP9O0RhccxHgKPWhYfC+1zmZC8//V3Rjw5NIt3lBh8B68zwInycZQNp1Is0NlhZSh0
r5jQudcmTIEhmoWtwGD/vaB410gTsnMCc7H3wUfBRjPbPK7ZZ94yTPjWJJ3c5bSSv2bFNnzFFLOf
Hwyux6Dbz98rqxydS70bEb5aXRjtnpaKeVA4i633fVz5/B/LhZ0q88p8cwXvJ+kLls1Svgb0PRbt
bSLFx0W+1YEb4ZrbyXTRY0RAPMDYnH2WmlnORT8ilmFYOFvZ//nEUVqbZ4K4X+njv0cpRqVpVYtH
Awal+MIHjP+sib2FUEp58F/LorwPfxuRD/I1NcyQiS5n6Blh+fRcGqn2WxQU7fTtYW4BoiO2D3z9
zl9ffo5Y+M5A9Rx5/r6HYs93Iyd0jQed72XJUDSt2ds2S75WeTFR/Vx2jAucUoni42xLO8aTuZVN
xg5GV7qYzRx7KsAjK1kYP49/cWJaAPu0oR2MBL5u6xH79Oj3EL1gW1wgkfNe+6qGL/kk6ZYGlYdU
byffopGuA5jn0Xv4V2VJdXKkB3dGYMjkce4cgHNgSR2EHHVpTZmwNcQkpDr3N2XzmceB9cLwL05p
Cf0g92V2THmubkPQDwSWt0h/ZPDsNxB8cQdL2ALaTrpuqMnVfrN9dmzbl0Hd4IhPypKqyaaYDdq0
9ceVZVqzt09pNJej3RaYPK0+DZVTUn/eZ9CxNv2F4VOxdPpguuxK6i++A5YjCgI5HT0lXz2XmxVO
WjOqNDdgkpFEsAtaqFDoon2u9UXIAaZf9Gd4+cnaP4/jjKYUPWBvwHUf8oFwVHh3tKDlfWehisDR
j7MMaLlg5P+YpRmlpX3ZKPQygx0DeuShhKEANzOVxz/hTUNsWmkZcoSC7z+aPH7s9ZRDlI5iuueN
R4dteZxyk5SbM1GLqHM7PSl8BMbSx1L0FD8vKHR5Qewk4CqVYMtIH/wWkJ0KpCpSr1z4Bsq7Fa0b
nY0WvRwUfNYvZ1HIRyaBDphVeOQXFvO5bx/JK5KVYfIcrdOnjNPwCGOwWTj+ar6xkVdd7PCxUjBu
oKhGA4FoOcmZRG0yxroSLDUDsTY0c8g4GqPNebbexfsfGgWOwKR/c9h9q1ra8kAXTENR+9naanJv
SsJNyVa8KbGpjjPcYhne1QkeatKOutjH6o8Wl3vNLw2u/sYw8+H1/OkrGvn1ksshggCLLHILXlSh
qJcxMZ84keQ0b5tbswKUFNLon9OHFVRVZVHngb0AtyyKQr+OREPI2typUit2FTSXQ+0knXNONiCi
oynY5OOR2dSjEszNqPKR/fOOufJRdSfzJ96dwN4M59tC4Gaequape5g7qd013Zxh/NJhHXTHeC30
iCKA9jIa9UnQO1+x5Rjt6NMUsStuAHD3ggm9qwaupkEfX7K7WqGpY9tbBGFh+ZOJrOIirHecNsWe
AGdLN9BqlKIDQxFZdvIcspQHMPCWBHkG+Pb0H8MzCl1+1gtTDJacJI3gycJjvesVCRHVoRgyTqvc
LM9Cw8MtzWu80riKxNAmdktPvzRKg2pafs97uhB4X4OXyu0ESxszmSoUkNC0Hregb6b1x9A6Sdcw
O26KxpO8pdHurpeNSBo/bHQ3nfXZS5ucg04D0wEJhYUHyH0RkEJTKg1Gf8DibS1dYncE82C/DZC4
N2zQsv93q49JJiZpQPLbTCob/8jr4qxwh8ayc07fcukFli2wbV67s3qC8UNreXNPWgCOZ2CbMKsm
369Ob3+Lgq6eWW+J5GbAn3++8KA3+fW9x7cvNMY7UEGvlClgW8Kf6RobnacE6Ut5JgTknnR4dpCA
UEyUWV0ySc3PkIDPM5utRokUqqreKjXfR1wIKVOPhTHUCn7FNrSjH2GYUj5fiKHIXghag8X9oCJJ
LdeOvYHAPZOx7a5A07EGjsmexDstFjWdb8gPgVDZkIIBkEUXwbIJ/c+pl6ai06HaWFq4XbyPzn1e
UsQzi18bkm76kzPy8NaBDr2/tP3qhZQorIq1dcPOb8g3RKaozfvsCZqeJnOE+KH7KcehCug+G4UD
uvsPUAbZdEFe2NOwR9jN6rWunUDbOQHhCFywvqDSOlOeuEoFPvU5x89v4vfe2DHbFtj2M1dZjPtK
APmDsIUEUlQQq/OEyykF+cXV0xWyfBx8BDRszHRVq/Ly5pNOfSL12/F/3tvD1bECu9W39AfOJgHm
wfxsygTu7beNMEp7fOXgctiTc0vuCjRz/KvRuY5WQOKQQGY7D9RnF8KMQbZ11I/ynZnnYxR1PDdB
0YcHOqKTUwX8aNPytPE4/JZ/IlhWKqYricnKo2e1PTFrskEAR/kT+qwEyHmO0a39covnX5YMcMDn
G+gESc6NBwEJNbsnz1bhrm1niLB9x+Ro2EW0r6DEKy2JHYXSptQWGVzl+Bbhh7CQYpITBaYQxa+G
XxuADx8YUmOdjmERfokxuSwYkdCiSj0XQB5IiHypxv6Zjh0Hw4PVTKSHtsyymb59q6u7OCz0+qrG
Y2jC+e1g591dzkCngbxRmiVUcwrZU/buzi3OMzZYeB1laEkMT37U/BBkXqg76eHIQ45fsysHdaKe
3he7qD3H8oNit4nAMjRT2dC4IwWWkPiYTiwEuIOVen6wgOLd1QaSwrdmZZjh1tf7rmltVSkuQDGF
Fobt0HIGmn5NnYrL0lm1pFxQAA4UQx1nb5u3/S+2Caf3ltfGY/A1BWZ/zspMHBwjh9EMwJdX9DeP
byzcgCqPphZjjvTD8y1gwcHE6w3Ka3UpSvYgxameY7IpN29QzLST4cyqGbgDpDQE48spKZlBWChh
/gn5tznttK00XdSKBkzKzqAlg76mGejG197240M2z4wXDRfXzHRNDZC401/3M/tLwJ9QrhX4dAMn
ztZuTgYj4A3RyQ0ApFH+SLY0EssYSG67xUNG8bZjQs0dyXtDJkfqXO5bEfEfakQ0BbCKX3X2n7+6
gJFmYVs7Nd2LVJY1CdEj3U6NFxome84cbagW7Fn5hnnRbFK6KDQOniY+6EgAfa/grtncxdQzbZ2F
aIMl9birehlJc67PjUmWPa29lsTtkbU7HNR310FFy8YG/wkjqOoh2xTZ0MlPhHVv2ZuU5ft+JGEp
csVupMBQcifnYYP45Rn8bXgCgNK1g6CD8qjl8DeBOppdso2hQLeWfpchg2MmfCsPEjv0EYQRhsFn
Ofl98bbbGrMr8nqFjO1lPiaLzooQCwPVOjpjWey3Oe1YUycEgPpwVpbGpdKz6apX32khRPfxHztB
YVYGKzko/UrqabQGu4cb0I6A+8O6iwkruGfKKWAOEIFIAp2Dd7rkP0Z7HrOrhXqPY/Df7KJ4V6db
QsP4oBKQ8B9+ysCq+Ukh6YVvs5r7M6vR4vPTwUgPJux5cfNUidTQJTtcwuKX+7alRH82V/YqUJem
5Oy+wsfXEnfKvF3egKgXzbBlbZJhRXVJ4/ezuggm3jpsWPOAKXi2Th0vQ8/nnCbZ8rgMeiEKWdIr
/0dQxhPvkkR2jwX7h3pXE5bfSkbUeP2dNgzeROd0tFtaD652dcd+k4ij9CGWS5dSzYXCrF3duviV
8uDc+/NUgTwHo3qI8+cj81mkFz6kXUqliq+aJYcV17QCNiD+gswaW/vOa44NZrP1zATV86ZcVNXK
5vMvO1eLMvkZABV/Gu0L9zf8Kwi7A8LMNoPUoLR8DeQJC5CIDmCf8Hd1cQS742nQKLAXZGCIP4+J
i4y8vujL9FRiz+OieOz1b/UYQxESN44qhNxbG5u8SRPRLfAwCB4zzuEPjPGDssXVobtX7tH+G3by
8rJSB3DLZcVAJ7GJkwDyR3iw0ZlrskL6nHHJPnWmTpoUIkQyAN6DwVeq5G2gShe8Mak5H3d1amrq
BTZbIc2hhjySHjU7+SzhGGbl7m568zmTuTXMKGK2wE7T23RAC6pGagj8WuzbUeiRL4E9hFxabcCa
udNdMW6CApenFQIEGWkVmKogOBWZbBceoonkQKlLxcGkFQZJuhNejJKAiDTvuBhnv2b1dvojPFnu
lw4884zvKFEm5fBdpHKyRJBidbDW+EJ1WEVetFQghAQUyr7vzDdfZk0qDkC5N0Wg1sWksBYi32hA
tcvbkMXplt7N+piV1jjaa46kjQKCPLs8KJmeIwejU5pakqQ/l3ngjgvtdZXLiixpYOWWoYZNcIIq
QCV9BhPc8NSP7Vzgr4E1gDNBdkm1akoKUDk19MvNYLRpFuCw38aSCrJDLO9+FlJcHdYGj8zw/Ipz
PP3YtdAad6bqjP6QqWr2pLy3SrItCglBPZHG3Sg5mX9nej/ieNk+xjgfwY0hWAWFE4oMCGHhgcm6
TaKnEdLLpcP6E4WdynN/crUOW4arBXduyKS/ZCyBP2rQ1/moOWALqCIM2ahAi35pXZOWHq5sgzX/
slQOxg0Nb+Fgz2hH17NFoHZ8ExDgvguikNdSEmrB1IhydoQrHvkjRv0PrwchKJcQfHIgFVBlK9b6
WqorF6JKCXIPMK9cZ+MmvXevoySUfzAXDn15U6SpElJwONaLjSU75cnYPrGkQUKMdZd8cb5GbtPj
BIdnYjfqkQftKfkI+JAQU+6JaXqWBhXxa1jsZu8J43jMn+7ZYWkYWqSxlnzPhY4lVlDF6ab6LHvA
4f++g0iHfXFmlZjv2yzOZmVIhThJuL4cNRHYT8g10+jFlKiNmc86mI4J9fbt+fc8gSP0gETeqoYm
GyJLl1wiw7g+DXRdzyzppos0Jd2KynIaX79UwSlo9SQK5/wosHmOh+MLOa7QuryoZfGNUxuSqOvX
6ig15cgPZxhXWqZ+o1OExEU+OVL+B0UzWT/svnE+cIzVmzh8u51XMjmaauGjwojOWMhLP9RbsrFN
tfjjQjTjJ7I/F6cmCDI+j4VIStlHKFnAHR/MaAizzJDeCU32WDLRvE66rUzsUUrjjTw2udHxG1GD
IfgLJbRit2e75Z36tDOePdal+R8/jCDkjQHVc73flS13WLuEDKkrdcmtoeJmv+VFX74qnKaWnk1T
BbgHeAnFW970xLVJgvTgYaYp/P4W7BGhUebuIU1x8tZGW92H7AbyAdnx+IBFSMKnbzL/rAfeu91B
Zs0vIm/e2w0LjjOLTKUMCOKd2fLFyJIwFWAkKIO1oRYGHCUr49fIWBRnUEc+TcSmFzBTqMXtQiki
kE+yAZ6ogl/khwiDi5N1c5oaOLkbktnWBF1/WEDZqWMUgzTFJuji/tb6IsTQPP1FKIRB907JDK0T
8MG5IGP2fmPa4Db+qNoFB7af1ooQd9DngV2+AMyqmwYJTFVhGlX620Q2UhkFyoHP9sDyA/2zeGtb
eVyhNt0wf2rBOsufdYLYkUdG5fJzFCBWlE0mGuClwjHJGe/UJtHCQVBk/rGGXWwhKR0B2UEc1n7H
Ej4qLvEDm3/e9mK6keKhTN8qIb+Ac7mwx+n6XYil2ADXgin3Jz7n/COTT96LJIFt+vuyMcpaoFpN
FR7JDDJ1X2SdgOU3JdFy+IrD361lUviyf5MiZm7lwdUZe+KfLMphAYFU2K2Y0TFX/OB11FasBNPN
9EiwtVslepNlOlyk0WzIIqEIhHMh2bwugyA4hUKEGTHChQsFvSgvK0tZKvkj6tScLTuA31HGl4xo
riAUfEdGkaTHKPjsg6IRwJC+8tj1FErO/jgE0GQ6eQiQRAvnmZ2mSdTD3QX0Qw5NN089unTpQJV/
XrB7wudBT6n+x6iRv9b7NbmRDR4MMvHYGNcHdds2aZSqKCcrBcyUFSptocxUFr0x0sA5b+oNLSRO
YJ0eE6hk8MCjNFEc7BU5qTZWulqPTz7NO2/Zee62oBsjEEKTZmEPnr1Yr/VHnUGH7PP4qSMY5agY
syTN5AGBGf1xaoRnJdpWHsS3xr/0aG/l+NUsKm7EPxBrHZxcczQ+pgJwS8j8L+6I6S7LoffADPR2
0DGLAH7kmp6TV8A/lgBFeyyfonlp9WFwswKrf8yptQGvVPAsEoLLQBNZ6eG0IAIYsrxwkTmAMfpd
2oNAYFjNNM3P+As1e77O22nMY5v5PI8qkzVsm80iU8F4xtf+PGgSZhkOrmOgngckJfTGjTKRhggF
WsUb4nEuRnFw7mctCbXgDubrdGLzkvojvrI/hUaqd4wTfFkgZPWle50y8Q0gSdPqfLURGppoMyZf
TdrmGV2aFVfozaf4GkJ1tlfGYDgGP+l2aL/beHaSQjc/LJdz8xz+Y6ipNEwEzSQn/pTdLtOx+Aga
9KKRmQ3yIld0SdGxXPh+xWjEQyGoyxmCb+/6jUZy2aP6Crwwb2SH9nYvrTOMegefvhAEM3N0qiTz
vP/w/womPC+Hi3wcwQh5Z/Q6QgmINxsSl5TcS/2N7I3keOPLxDQoH5h72oCM/RqCCQH6eZ08zwIc
OA5zdvWiodvaPziEs+WlRj8qO51TkLyx9yoNMS8M0VPsQpT+Ha5ZTf92vlXoaVVoMnkpGw6K2Rzl
aTB2GX5HMFlkRU3LrNvu9UhoF0WgX15h70Y49vzwKW/kJSGdeRoEyvRtNhkkh4J4gf9hXIc1eqUI
ZavFfTfWwv1pMWzU3PS/Vf+QnQzi0tWM6Qd9khLpDISazkLkMX9DHovnM9O3EW3F62T5YJqsBaXu
KuvvujkFuw27Of+bS8exuoZfhzD9BuA86Bhh2Qi/N70ZEJg+fkon4BjDGn+Ua8ECii/7Gi49Bw4n
T67AnqxYKWTgLQzorQHPG0nxS22R+L9RVe+y0gD61mND49MyJV0dS+rlawzecPgJifx+XvlcvjQP
XdnBfjJrMkGwDZNbnVUgAeM7GCzZaeaSMnQMaC4Wviih6iNVfhlRkDzfAitqxiSl/ZJcnFWncx+Z
uvgdEea5CoFR9kT8JCTJGmUSER70hnsGsjstPOH9vMCOBbMDcSb4UUPYdJ2QESXdVfGzAlS+4SOo
qq3oJLJ/QFstGzVPwrzfaX78NN22+IbDZ28UGF3zOJ/XsahNTWeMI/SzoT7FSpLdA9o7FT317OfF
3nZBVfsUuFIaXPXNzfRuOm9LYTM2AyOkQCvMbZJoN8R1n4oNLfkwA1e3ZtH9JNqJ4+rJqW+LFBSe
M8YYneWlz5dZ8seCELNdmBYYKpxOPvsz7LRo4S20V8A+ake7G+KiEEdmvFp465H8BjuVd95lmq5V
PS2XkeUymBOPFlS36z84EZKHu8f3jhZCh4PttDtKiZVc03taOzSJFgI597m4zOYn0F0pMpz6KRMP
7i1uMiyWgA0S/3Kld5mnPe4tjBLyqObkXH/JJIj1iPxZWfkv8KpsgqY7X0RnowQfkBN1lZ+roMDc
w0W3qSAHBDkK/WrmDa1x4K709awMzAUf3ehyH4JXhd2jqGZ9NBa5N6iMBfw9eOHH/fcw6D2WOWnG
qtRJoUXzsNEvC5QOcJqN5X6XcTK9Fh+5RBJKahmiz3KYv4MFXx9zWYZ6Wjsqp773lY47GDitdIE0
7BNA+fliqOB3yV9NwiG5IVkGxFz0QE4le9n9NACGn34Zfp12C3zxAp+1WTPeXUoYixT0NOlBMNgG
xqXGQcvW9t8yewbTj2Q+sC61FdJTAW0Bi0bnfti8cd9VbhITgaj+QuFFZ0VIfDsu8vp8EhLjdh8y
tVmrVsXGn9ay7xF+ECWzN6DpIDuhl3yc7h8FS7czII0Fl5ivgHBmWyBl8PJCXWbdCXRrEYrfDO5t
1OH/uV4jG5jVdQV2uS8AH3Mlg97+b7vJAm1036qkEU4LMreby6o9VBNdKgYKPoASapzDzpwGqYEJ
4b1LkNl2y0IUtjeHKegfJGVCE34wGCLioEew0+IOMNOpXjEwWWEf+DnHxAtWFk1LVlWyqbB2AGck
NNMUulqM81HcDODDLwGPwNzYe0v1a3s1CZNrSEEJFk7QKV7U3nlp7kijhiRZXbyaP8mK98Rz2bvB
rEx2/fN5NkNk6A/TDMKZgMSqSeTFhXKdTTe9UebrtdV7YoWoJQgBAhpIekFdx9q3zVJJSUbc69Bh
s+DKHy9SqyFSb4+nEy1jwOLGbG6BtuxcNDT5JoJF0ka/G8VbiF4PD5kxZYsiIEEXP1EG/pTDABy6
PKhGRY8jLMIGbUxOjNbvYM+m/EbIf8SgbkM8BJis2e496S9XX2Oed1Rdjn/CYLPC7qh4zBat1DNo
67FDS/nEvu+kAWT1eNx/0FohabYMjhqojwPA9eJGU6+AOWrI2RQ2659oUal6qpd/iLnjHqF+0WP4
K7szYJzVTwBEGHT/6eolZDECwXKMmAp5/88gtecxSx5NTkHLFa7ggF6lVYUkZxNSrBYd/9FnoGU9
58AIRFBFtQPI7a9x8kCb/WHJDDA+mGzOBnglHHsBOleACrs71zbHngKPaR7PzQMIVRvC/p0cobSt
BC3gAKB23/Ky708N6f2tpNuftwQ6Lq1mu4CpEJO+9+ehih0QitPTVoTj5TEaPWxrbIXMuFXex3pJ
dxoXyMBJ0DjRX1ryQ5YAjdkHwwmUG0tN8h+jKj02v24XHJxW2wwQvWFIhexlPbg9hP0/Upgb4KAN
tc27EXiOsfI/54d0j2hUcX8+j8ES7AmyFogJD3B7/L5NjnkATYs7CmDQ9tmStBpjS8m3ph0tFymN
AqP0Wy+faGihvAGFl22VPw8cUYwhqTxJX67FxnXn8FyD9bYksnqagEkQsvlz8XGJWucJZQLlW7fE
7KxjgWDOTHqgurAbtBaA38iNpGw4vfk21Gp6MJq3hL/6ReE3jxlwfMy982Nxm2UcgbynRL8WOGvn
rIEJnOyJvnjDvAz/hn76ftmVPPF6mTUkUNDsf3E1tkbPc28+G1+lah/KCdWGkgfh4fQMncXmCdlR
WFE2SzVnG5ry/opBqUfVrk1pSGYOPRJJw1HrQysFxS72A53rAaonhK40mxWOhAtw5ZBjSrZCLlFk
nXXoYs3U0Tm+4wZGp4duwYS75o8D8+K8yF2PXgpwQ97ZcvmUlEGTs6doS5Wq0nUcDg2/U46XfQfc
vsTuJe/aAoD3MhzYb6V7cJaPYlNUIGRUKGiZhSmxqzhS+cGeKjFfJ9fAKsDI9kZgEq63Y/y/HT0K
3v9UM7Z65U540xBGGpCATwjju2SKGW3wjeVt3/EeA36NqysX+irwutwP6Xh5R4VAyppMx80Ag1Ny
dO+zcnCg5vzU+qfIppk8tAE3l9RGF9sEJ2c9t+67fY2moPTPE5jHWyi7N05QPSm9ZtGj9AN/8Wau
I3H7n0JppPWRZ/1VHj49tyUoeQufHCiRn/L0vkriwb2PESikW+o91jnhKEVsnmIUdth3q6w+9m/A
5e44h8pADMz9BfQFhAfy+DC4UDlKWZEdWgUOU1u4WpeLcM+p2eZKRLPvcc3LXiLg6HafukJW9xfA
NbxgPutz+A/ojVtU86W4n7Dd/catW0RsHeNauiFSBmwXUg6cfV/fqQazkXKjWByzC4yn47dNIGmr
OiUijiE+/DJQ6eYhmXv68w10M+hIfQnYBMxjEFZ26qSnV2b2dI8+Gk6DXD5ZYqZtq9SfBhHMmGPW
t+pMbQ9Yqgi/EKglDW4sgrVXZetyYxM6jhK6CEj0uJM3ZsYg0I0EzYaA4hwT56flyAn3NR/MvU5k
A2Jy88AgvCcOCwqwYk+9/U9fOCQCsZWLPxean/w57E0/iV6HYhT6KObt7MARLovEUgeNVo1fhzT4
fjTKHQmWQj5tWU26Mz7c2pp/bplMdruQwRniv1GaOkOIqoU4byOeUky8a9tly/y9/QMaYQn4Tfy8
bhDywNVL1bIopSA1wpV5rOJpsHhZEKtsgQVwqc0tf0OL1cj4k0nZsbdOMhfsfDya9uPoASg5focl
MZFROK3pIdP1p/WNZTs2oykqvI0nt2f+vDorkjHloKV/SnCk7r1iXRw464EWKpfYp61RQmdrVDWi
2HES9JU5s4ozoMpwq94s/IE27heCv1lNnawptQpns4Sr69YHIS0qaDagWIy3vMfr6fwmrFFiEgor
Ozh7AdPlIuuIzxYH/3G/QL7Q4I72LbeCXYwPHowKp2UMhjaL8EydcIQFHtvBXK1T3cpg8QNJrLv5
vjnSB76ciEopXhdswdyyyD9WKS9j4lJHMHPDsk8G7jSQTCyHpT4/PuH8G2cPw+/0qBeCnQNZVgkU
FpmDP4eP/G65se2OllLgtS33jex3qfg9EMmJJF2ULLBYZNwhm0tvzhAZUZzFC6T7u/XLEBnFkqaD
HncCiQ2EsBAq9ym958IQHyL/WZOJ7Uvf4KP5/J7g3UPhac/2NPHON98rT/BvGleAzYrs2tZiXEyx
KhtRRarph/OHR1d0eclkwRP4t/bV4jtwvDgABmM+iLEX4mV9NhC7NdXfnHxygiiepyMB6dAY81Gn
9Hjdj7cFDPz8OsD8f9CCS7t+KbO1D5Xyk/Hr6rOipDL2+rz+sFgzh1Q5VRcx/YUAAC+S1Dkab6q8
+T7HDhw4Vt0cnIzAVTHsn1vsf9EPnrxfr8CTwuDwNSTqZ57hh8ZQq+eSeudlfsKOIpolHlnkt3GN
FZwrY2OH57KiLmMBPa9OpjCAKJUB7IlMwxyekVJ8iGmqIaz3NqZDcv11rr+6Nhjn3W166R2Pmkie
tuJtWrnFe9deMpqgT7O44sM65fHH1RjNdf0KYG7yTud2209zWnss7fEK+RE9zob0/A0lEdzUiPJo
Sv3wHFNwEwm4koKovPGY6NASJhpzSTBJSVCs6c8jIHJ1e7lPUejpaq8wEYsb9hJO9SNW4ozA7OPD
VQjujXR0KDJXQGYcbZSVBXrSKZHUpcBWUXfyODI9dh5NrJ7BnsD6u/umdSqChkVhXZRNlftIjSLO
ub5TxnysLSC8TnvzDAYV5CV4+NIKShUum4zrziCIYM0b5kv2tI1E9JC6rAe2UaX0IyveKYadCoVR
s4i1y+0uC8J5m4MOAcjfTmcc3MU2H1//zNfAN6yl8YD4Ggd+F/GBcxHNhZNoBQz0w9gNKDvLM3tX
8jRq33ZjXi/g4FcAqhHxvaEmpOs7KKyylAiyNAp2y/epVmpumc8esudjI/cykY5L3Vzk9JM6HdKh
BmOPoVGg2UgtSJv0PH30M6QD04iXD+6gaxcRsNZL4ijSDGHQdfCWReygIYTkK87zP/u+lYoisvPu
PRO8N0lVC19FNaKbImzALVlYC7L+aYBtgMwdaDOmYSZ7aEjiF/w3MILZDhG+fUJxquqkKm1kwhqM
QMq7x/Nxi8WofXp9u8Sn5dtqOQCAWcf7pREiPnsVhWQ/+TuIZ96zpqujucHx7b/grTbnQUi1uG1a
+It1TcBwlVFRQqtvU4fexdmnWFZ9T3DK93RQWgZrmm0SuHD+0zVR/NkYIIAasSwcJxNSXVqCX+W+
YI8EbUFoB8YDicfWF1ajROD3OrLfghyjk5xcwb+ZTcE2EHQTIM55RTQJyPexUBrDrpw/CvsMbbTd
eucaRGpfH70VmVAM8yLoO/+165mma/XnPNXVhlqCWaLpFNJs5CFP3GYHvvi+4If2Uh9UeRaYCaoY
kLpcoSwsJ+saUhrXETgiDfnYzghi3EI5bRNmd1VG2yo0RKXivgNlMpyMOnhvobVo4rQSQorw0mTp
RYIHIsk4aYaSnmgZ7nDIDxn8s1zmE8XREfy7hPfB1CqC7mEbHeIX/8wxcQ7slc5r4WGp5aEAHPd4
Tbbvkjk6U4+28Frwpo8KdTGo7vWeJTpJ/401//JztD8DyPP35XoK2p7FrWqL8JP1SZboRtrKnWzM
zzpj+0RTllpjBIo4vuRh0ByZaWcEPmkg1eP0Rrx01F9W8P8OQZcLquCGkWi3WqurhCby0JKVq4Dq
a+cZFWCXfD7thPyLK1ITi1k9G1LooygIb/+O3LFbxMLYjvFr8zl+iRLwnxPhSBOPHYgPpF4h7Er5
2dBXA/ioW19YhwravFN5sNfXpk+f45zx/MNorl92tiJyQX/DTiApUE96sdhn2Bx22Txm6JjxkF1a
qh4X3QGU8nQeVUV45OnT7iMMERMtdNX6yjguYJz2xlYNpLaOwJLyJun4sFraXNBgJ7dd+HtPn/cd
evsuhyNxqKB9JuXbj40uW0xanVK2GFaqTlq4aYq04HjpkumM7GwJt+56z/JLlyRRQ3JYfKmwWX71
l7QHGFs11X+/mnzKCWFtbK28CFWk9trL7rw+8IdMn4RXL9cxoU0bROY1nT63mm/mAq7GU0nICq3X
UZKI2AlNO+dLEdCymNWaK7YhVMjb4/QD0DaR4zu5kzydnQH+a5G0BmBv591R69A0jNZoUfrz3J20
/DoAiqpKI5w+zFEJj+hZnzV/9eH74KHD4s0u8P97gkzkI8NbXj6lpmpzD3SyCelkgLyjJyqmlBOD
Zl2/fLuTboiSb9+hPMgl19r7Hc5vfgt9OF2CaMyd+GzQw4fvj6cuzlMwmNYLwR4HZ5ccsIT09ypj
8HnmdxPEEomzvq1uDBZn2+CKOeXSYjDcJG9WuxTUQbYKXWpgaH7qUBJtfnJ85WLPvf4lYdQZ/yDy
6vCFCH7cj/vD5HVWNFw/lYbl7EXriAJogBKSnTrN5vz4tdTeB0TtwJZRi0DRb8yDAVNNI6Ee5qQL
WcA/jKG/B1BovhIxFm9g3s/KKS3i0VhauGlgK4yfVuFL3op1dKMSFneg6CdgO62JLe9X5wEs2AMI
KiUgAAuwfl+WaYWGNzZnLAd7hflZpkrN9W1Tg61ig170+NAbU5bCwdcrBuTDs1aoj6dt4T+Thus6
1WhaswY24/mysmQyJBQLgjW/yh22SSkCVO6opReQjUODVXLkkH+cxw+e8ZMYNcDuoZfApOincLTa
R2ZiI6VYuzGj+pJqQZ5oFI4WAxGRp/yYw1xhKeeVHJAX+XF/rV3MeheKRe021bgH/gwAErKvPA43
DiYsk3pvKqJM5sEtQJVo2jkbg6jj8MoMy6V8GWbtrNX0JguG7ZyMWGpO7joyFb28iGWpNo9HC8y9
UrohvcD0xGyylq98nipaigHTzGl3fVykVEtR8Q3x/merYHvL0NF/BNec5NuF1Jzcp3r7mUTVNwHw
E0yq0BR2d5C04aLRQ4/nQAxTiRzAxGcyqmdsDZly6DJyOLK83D2vy2jzWLfJzVKaKVJK7ik8QzV7
KBV8EO2fphSpYwBdGBI86LmDJ4nuMAAPKBL5NhX9I4vNundz5eY7WevLbzbCkm69Ji2JydC5z3Lr
C1klOQGGiSJowazvLYFGfhsb85LKUG+Rn3gRC23wCoL4PnWoV9LEERyl821aTzYJmjgXbMuDnIIL
MuQUyUovy++/M1HV5rCumCBgVNbOK4Yn7ADFn2bU/n37OW1jiKdauPBJzn9Ok3V04d7jG/lOCg0C
ibmaE+HvdQSKYXISDKGXFMOv6tAE/oqNR13BQhmP+0uYI6CYjKEOt4f0JdHjdSXzPLct8PaNm+sU
JkRbXV2bVaH6n/sZZv8dAGrV4ZDkwzgJ5ciYWW/1auu8zjw2up4gX+spkFgXh87B+yUasJznmPLB
aCgL0vs2eytv2NYKhiZrRLPzKE322pEN0ZD+0MBsEgla1R7SU1QjDed+EuXpzHlc0y3HugdIqK3q
C+mtUxCYkpIB+I6YNaq4LbM2Hg+nKHtwwpGlbUlvq7Uyn5ZWHgLr9cbF7zKkONQf4gW8wiXu3JDZ
09vzPTUHepl+OHZ2cZrALR0vtmAE0mMYQ7VW6BkCCtrDOKGhJB7svPua9CwrCRd6knFg4Q7agmcW
rVlIKZK6wcPUqSidrybN+qbEggy4DidF4boil1TZPGq1+6zdVtB7vGuCml3xzbnLQ1w+xYXszePt
nUeSwAvXyrf8Fd0Ll4zboVqFEhBCXvxC1O1wL/aHnucJz98y5zoXptDkzCNlICpeL+aVDSvcz2pD
sbVbat5SHsgvZAsiqPtKQAasNgzsriI4xo3up3oG3AK8N62REE6nV8qzZcaUN3KOZpMd5QbBQNXb
7Bh2If5RmH5KHG1KUx3dY60bGtLBRXWeHa1SOXOwWbnlwbqzbGsnWYUJVmE5hFPqQXA6SC/TPdN4
q2FAkVjYxZ5VNvjTMP7GjdgHKyIPwuwWDE40PEiBjP1W1+e1BPYs2c13pnA8x4dMNx2IO4I1KeGi
gCVPGkg1eRxAvyLFuMY/Gtllhpu+AsYsNhWcap7N3gKzCkGL8lVxSoFdGX/gXH345K1C52q6YlEE
kVEyVm1MA4J//GFrmZw84mUflNMALCqtEfwE2WPy9XKvd/4HU42l/eZceptkqnWoZmammFE+k7iT
gd2IV7kZkc/95tp3yFDvBdmrroT4InlREjFKZxfLEd0yhRPlNgMyBPN+7hz49Lu3SdXfnloDU9uV
opw7zT5rhp8GdyX6QDd1l4+poNk30pNIsRR6cokvY869A2qkOftXZIt3mjcd9vGPfKE+7z3vd6o4
0g61FoWyshu80GZpikF7r1bC2tvntMlI4XvFnj9oxty6kHzNh0pnMoP2dgWx4RyyK19kmPmf7G5p
Xfun3SOeXSHkW5AkTN3vYhdAuUakYs/t/pzoAieGcUdrfTOsUf07ottsGCKtdugMQpK4XGe1vydr
lafgSjyeN4EuHiwPb05HCtyUsnJaFzrxbfjTLnyQpNglIAXIgEhLePvlYbtjJPjySl8fA25jxxSi
V+FfF6V1VlDD21flf5C/Ugh06ln99NuhNC4Dc4l2iHY5CuQQAoUQe4/S5alawTRMxkkfN95YIOJi
n4hC0Nr+0yOql9x3YX1EnSR/qxtjRvxojjedRoQ4uUysjf75LaCAM1o1ZDe2Cm3zN8J/tZb7qeRC
yqaZBnRre6LsX5SPiu5X6/93B/DiFzYkM8p703Z6bK1b5VazDvocgFsbPs9b7Q3ejxh5Uax+xxNz
64W8uysgRrtPJGunHT8zB+jLlq6dX5L2L/sd8EbYOPsnDZpXuDPcx11+pL92tphUb59BoG0YINg2
gBEBlVstdy6xuXana79iNy1RlKcy0oVCIkxx5fjtEg5AEUYxm8ksoBtGnctOf1hk1MJOmCLdH5pd
vPXRdfGmKGaRc4bcyjYAQhOO3sqof9P2pk061DpAxztXbIIvQHrjoG9BA52baEl+dBT6ChdL/DP3
iVJqrfKHUlxP1EgzUU6u4MupEKO/8xMhQhARXrMydjwN3xGEZWem++LXzUkD4q+TfaqPqdd11KEx
XEITw1NwUBjaFKfzmtawiSPbspDRbcya/eYSS6XlkYK9rrW3uFjVNZEjTpoK2FzzmMph3+jzd5Sb
H9MvAVef3cN0QitHq2/Q7PaQSMwBL4BshYRMUfzy7MexlNdDE/AFWvhJns2xdRTX3mRcsx2gnFGs
P/kf7YkyGAJxZ5IT8y8Z3zJitl1w/PposTYZ7L2V0IotjkJ1YymzgSyxBj+AmzfNUNedz8oY2pxp
iuVTWmApFGEAEN2Dlz/LYKrdN/Zlz/0gGExINMLXH9O9jKqy2mQVJ+ITqS4EjnlEhDk8PJch+XuV
zsLiEWzGvIU5r0+h8Y+7z7lNankW063ULzU3xqqOd3ImJV1nz/nkyN42BJC7uOXyzoTkWj+cDbq5
wk2HatqVIpe9Etd/5tbZrb/rsdgrMNPxf3fuxn33Q47rmBSbahV/95h08oL/fG8/YTcWN2OhAEB4
uhxxx3hpTG7gTCLIL+a630smxFZAwE/bEaLoGvmba0KwlVq+As2Noh5coPVZkdJLGyLoNVjujwyB
KmT9JZ9570w1bJyB7yEmWq0ApCvaHe8sqigQ7SoHYCUMVwif3rhhJtqyzFPNhXGDuOVqiz3L7xV7
VeF0BAxl2H3kqNsrvSN++eUXwMcwU1v2O8MLuUcXXIRg85BciFw9oz/N96m6ebxpAdgxM1meXUOx
Iz/CR5mRMOSNoDOY+3pInkr08aYuvYdTIb5JDyuG0GHw1rox9yeVQm9t/EQtOBi2K8sq3yX6tIy/
f60SG5Q5wZoMX7mZrG4JoM97zRYih7Z4/j+G4FOFOf/I/O/DfbfYnwM+vhj0urJxoRkNaF6Pqj7/
lJM4yxDqAGeSpRb2ThLpECZ34aB+AGVXR1tcpKIcF5LoN+CN6Vy1sCBPYoQqucatCC9xpzupcsAn
ASqn3vla6ySZffwCV0gSO8iom0R4DJdPYg2LtrT/JX8sMNNwPVWI5ZFGUCuaku1hHfiI1E3NtpQI
XGayuN4A2zYqJ0owEHj7k/vpQkzEkCgE4kZuJAqcZ3QVPrk78mZOn/uVDsOknKKK5Ndob0HdfIji
VocO6LA40jngoR8HEchR2I+61bhCUeyefqha3MCTQoAAoL0uXQn5O9m9pWwfdbENoPJsaQE8cuE1
WA8KVT2AiRqZ2RYYsWkwwGVYz4ThG/qeXbZC0r3RwlKxfdcYvBrl5bILTb7utWXBtNiDeIGQmyIJ
OzRoWTCh8+bbIMH0DFow0g6DWjz2g3T6RR5Ueyi+oYMCG7CTpyfrrQGifOZx9F6oeQP2I8mSew5w
HHWNRZJQe8sFctqdG4mxN4Tnn4PCtNxfrESadMcP7Z1h7IUEM8O5AKKnUDWPCDsTlSs7zDsiZQaO
QQl6vCbPQ939lZdxzgJo7s0ZyJUthBPkV4mdffWhVBL1/K9og7F9G3a5xpEunmxLm/D/p08JJ1HI
Ogd4SfE7jsoD+4sBFKVAEitUtZZQ0Tp89lnLVWuk4EG1Z+B5DU2Bd+4k0XPbXkhEoYzYzCw90JKs
P3vnL3om3yqwU1veKP4MffvoahvaU9qJzGzHZW3FOBfZfgZoLMAWGqwAxH47LYFXVkDnDkx382Cq
n9BiUokhtwIin452uvggtbt8ysihWgE3Lf5BFRHUUzySCUS1VPUR5LSTwOio44r16KBmNIIeIl0o
SJYHa8b+sHjdxKHGqak60dLlUL9Dt5Mefp/q/EMUsCPIbUnavjSpS/fh4OVCYieCuu7JfQ2dMdCE
rCTxkE8Tv/8kq0dYwkA2qIIbGleOAqSqAKgDFYi91d9iXwvjxVwBCLfCxb30/Vw+LBS+CBTNVulD
FwkVeWoywwIKV9dvkhlov/HQf4E6HvjNr3sX0nxFqktnWsPEwko5vezlylGBcGGbgbSNklduXLKe
oz9TD4fplCsnuxVWjo0PlLxTTdq/AShlJmv1oKJkxBds9Sioj5Qr1FMK3TpNrDHbwqR0JxcRXAPA
X7g/9oOCE1m2tgSuawFd1vi+uBJwg4M3ET6GBgxLYMfXDA4hH36DuD+nSm/eBmluFDOy+p1Kwlm8
RXqKhIQV+lHfYYj8HFxHOOsS8v+34VvUaIrsLcig6DmfzEHJV71Idd57uFZNFkQcrXwNn5Gp+8s6
t/n8AnnOMWdXEWvFZ14KBK6mRSfPC5055V9NIYIRhdMQGxWIDsqhM0Zm1Ng2olNmO4Y6l3tQMBlz
k+33rdimj1NvDt4Ah/kEil5uqiMDPKakOvK01vdH1IIaAX50/TtzVOAS9nzrqCQzVDXFwaZ2H89x
942+VKuJyLFNjq/H/pFrD/2VLYJQtwEP0a7Aw/OGbZFB11nsQH2uZHoOTp9ygN0vD5GW1+xbKIcL
Emo9kgkOVHRSnKRpGJcidGpcr3hx27YYziECVFyDnl+MqsxjHner4+dnA6cRZDS9iw76pxeDWUX9
IxqWaTGKpRtNMyRJoOp2Df8uqIOGVtZNT5/E+CGYU9D6oVcT6HOZJ9yRs+hFog3uGY6TLxmpsWJO
ETnGOsa9LhBNRuxLLiiaSbvf8s//vlQnPsVGiLTyYctYWeRKV4bsZjtrQf6uldGkP7RuM9V/atvZ
0DdqYLFU0O6ZZZDo8PDIUH5O3jltt7VN8jOhR6Fvov7ogL4af0tlLBA1I6oOseozwaHElX7DP+8f
BlbeO/0RhdTRhc8puA6Kuem9Xbp9nLw92syI9DIYPqVjo29p73VZ9dMe7HBfRaWiAoQCV8Iu48zs
HMri/XLs1feYButzK5MEAQAbQG08ZFrdcNqGhiV7FPFYlnwwTdDEO9FhN/gQdc+vaUQfO1qpmng+
fq3GBeFBXNQBR9VF/hJ17NDA6PZRdari4ybE0XxmnOjgBGx3oSheLaJmd+CcpabFxOvyqO2+RW7w
V506f7uh7jpeYist2kD9SN3DkcrrjcGIZ3qlPBYR3odz0JcYT2L/PUJ1hSGMsbxfq8t9au//Wqix
JR4xKOLO8AhkomrsiOHaxrLKqRRJv9NHb84q+iiJwipH3bL98HNf3iqh+d18LtT0+wio1WQk6cXJ
RwNY7hK7sXXemafYH59L5fT2EnCpqFkmpiJGok4SUajeDiIy37TuYqRJ3imIz97aNPi/0Z4udyEc
xxsIlNLXxF/8pNWOD+Nbv5vFyGFogOY1GBm8cJr1qLNKSI5MT1OElGlJQPuOfbFbOzsjVvuap4Gl
zO6HkjdF6xlT9dpEzWasQ1NqKy0gvgVMrE3oMoJDMbgmorhzdoYgl6oC8bduC8QxRw+XumbeCXYx
1Fk+hinnHJwsIG9+hJOyRh4PKi1wAparzj7d54xRx/IDKPyNWHeBzdn14qLluKrfcK0kYIv38s3J
CEucrIxcy5wYGnO+2tRm8+U1iH6zJ9BH2v96BPGnnl9rmbX/wZbyxI4noQt88UaVAAYQj/oBtdmB
ApJ7YDPGgN5b7bCW+mAOurgSCkb7x2mkQmGriYhfsj1MmZUvT524rXgvRU2Hp8MNnI+8sSIsLuPH
SiYup6j+Gn9Iu0XK18OVvmJoqpj2OInCAcZiq5WwG75PtyAf6Gxcm0LQDY4c+v2kuXcArGDrwKJh
FdIlsjPVI3tx7XL0GX6IRYqZCmphlmQBSd/ZRQM+tRMx81NUaiE5Px28tKR2P7013am3jCeOA4LO
ptzfKeJAgqLg0W4xNf0H/VcU1Z/jdYu+qSQ+MtYZ7ejxdDxVOkSIHidnJajXOKzW9jZ3QaSb++VY
9OHwBUyZZCM0KAfWUvtxSSlQRqDzHXoX66L25wHlDuj6Gvtfb8kVUfTMl9xaCb30KwgXksttM0dW
3MJaIAYVfUmMbsCq8mG8zMTAItHPeqUNh4zXrjuzvW0RCQBkWEiJVr799XOOBYZEUhZwvEWjCynS
Zl58L6eYDio9qU0HI2zz+yp4QufF4KC0Ch1lnC/g7YNcVhotKfBYiHUNVYu4iBmSwEbW9RHZEuDn
0TnAWx13klna+LOuBs0AkJ5vIYtlVkoPxfGOfp3q0V7bkpD10vcXqio/GTUlrlog6KLLROM1sRYR
LhIPlkpCJTRV9ihFHi2o9wFXwTGS9b3PaxDLqKlUA/WlhaayMZ5ieL6S/19TluMVrPFSlzkEQNal
8qEMWV2B/SlZpfJquGPs35O+21YDPsxjwul3CQaEkBF36JAua8gT1PzPyRd9mpXHr5aJk1WIPFT2
tH4KLdMzwwT7JzTpv9XhwDxP9aN+oIso5o+w/H9HZr1joSG+XrNxr3KRDfdTOHu4lyDskkl8E1/s
lnnirzBXxbqXVhAzUKYjOLKRn+xVzY8sSU61S7BoECNA8tAibG+rl8ukdzvh6urJjuyzBFgGndxd
ll1EQdl5EuKIt/scAnH/DyEBmocQi9Q6aKIt4DDXqFbqHSvpWackewEDbrninVNzMCjkbvrV5bEE
/e25gLGfTSUYtoGpn+D4f2jwIznx70cerDL2aLbMyBGk0nuM9D/Kg/kFwjjSHJQqJehvskHToNPc
6UVGAtfbtHIbjDO8Uuq1CCtN+v32WVrvd/YZUSkNn2J62uYyAzTknWPVvmFUbF8fLyaEl9F5DExi
qaIhJDD+WlohZuzUSYJ+p6WzgVtnMeuWvv3J/ZzdLIEmBhb7NUHPNiKhgX2VCSczgaA1SUvZABVn
cA05plxXoFvYmXZL9M15JzwLE1ALnH1hl2QP6wYGrtUmXKjo2tstDmSHt7l9YnhFNuzsLZmIw66w
fuW6CxIBQTGZAyk6a4/uh7he3JIYu++d66FQIU3MY2ORWwy/qX6oTVu7xNhQAoAlUymsGO1P2a2/
ldNo8CZkgUHZ31vF4g2DGgtFYfqk7Lt76HS+suhtYQdEjMegmN57vjlCHogKWvmM3bxSf6fq6bBi
GKaRhSsm5SP7R0bvy6DXSA4p4blHeLOC09Qy1705GJo7pN0x79WTsaxNz3w13/ld7tLrUwvKPYNW
k7RThq1JkuV8eUUIG9qK+5w5PPWZP/gB6RahgwlTRs6cIhw5ZL0UkXDPOWOKy3V33yDP2roxxDD7
quxVCuuOXtbulT0B5C0zxNBzudPwuGu8UdKJ1uA4lqgaH1Uq6UXfIbIAE6sUIZYfaBDM0cSWJH/h
+O8ontw+d2i3BF5RhBYgWckhz581sbIIBMqXZJvgYeXQW+8/oXwv6tfWWsL1EhndhMMHA377rHSJ
T2QlvVhgdbwC5B5o6oLLjIMDMERqyPQqPpss2IppeZwZQ66hv8HTS9LRVBhhAUjvJLeddRev1yWo
bIgplYlVvg22fpw/z/t1LCBvvVqcCeR+892Pl/8xoBH+mo9sS4pYgyUFBKnXt/R5MoE8ljthpgCu
h5I7QJClaxP6qiwPXILYkyZKPGB8bQ+UIbAKgNOOloMIM/zql1ApdzLy62Hr/cifIkRKAvIhHd3d
1o1Bf1RS7hEIKSTA9oZByL65hawNddcMKdvCJPNjPstazRozs52XrD19udptbdaNWdCs04L2qZDO
uO/wO2LiMsz6GzzGvKj8GCO1enSoZGxHcOdCq7NdlZniApsXf9ltYhYJWapVPbR5gW/UA7pnrHwf
LhPieFwy8Gn1ssJXfp91G6ZVolM+vAZ1Q7FMzQJQK6YmM15+WS/RD/hV/OQs5aScWa71eMNSPxGR
jGQJ6dEaQQox2Xf2g65CUpg3UzOXNIP7qYEL49PBbsdMHFBHxfrbefwU0v819SXLJy1Kkh7kRrsI
NqGYC090maAn6HlNUoG2mSkPrPuvf2atObVO2LR66W5wcKcq9xx9jUFFyDKuTDa4JNl0yeuOJZNM
6BP/lOyDaoLN6YWc+DPuUGDdsObKYaENnHqqskabU5gXk+Ntcbz2crlxmeYVCBJaUaTAYBORPMuZ
qN1Xd9zMy4BErrEH77zc5rDZvrjyTc7QnRzfPxPrhXwecoVVHGfIqHq6P+4T5RunlVdTjkuGpqWI
SGw849Mu+jw0FojXzll/lQfNtxLwBVSSfaMksfZ5A9j+7YQyTugqeKLs7KIhYKBp+N9kA2MMEUWo
q5eHwzu2TKs09mqrp3UKRBDOsn2yV0R/W3uFkNRpo2pO/RvSDQ/8LIvQQs2jSSTog7Y9bH4DnQZ0
F52Kbh8NXoIRPtK7WfEz51+1tRn6jPIjGC5SSW66rq3xyk+LIQEtFApwhMwR7qbKwfXVFZjqWA89
GodqeoGB8vTiGlmNhryMiFA7wgJHEh3/2qbK3tcXd4arH2RNip+h5XRuVDW711V3jDlVj7Rv+5MU
Vl3N1CICi168mcgIt+QKU6pjaOxfJEuFQBBk9w/Ki68cf9BMkpHdm+siGa5g++VHgop6n7yBDR+j
cv18b+Jt5R9KFEP7qFx46ELHzBDkbfsZLcLZIoiT3tBnSqAtsgHIgt592NAxCCQaTFtTv5qdrMlo
JoIm2DLkPri2n/MXuHfT0R8HhIMGZMiIgzjaRmCL/i97HD+lXqbfHQoaDZUt3r8yRpMvMYKmKbGp
1aPb6+jo9Lgj7JxURT6/cA5Oxr5Wp3NWSKHZp7PLqwT7CNS+c9MaPE9jXBOKS6dZAp08Ek+8l0QN
Oy1m0tCCSc01L4qq1vV9Olo7ssFlT9ZVtN42AXG0x9NVqYHYQXR712+XwicsospyyjvH2SLlwImr
tRtAQMycJd4Wz6Hfyxb0wadLUwExWyWhhVIU6yXwu8p0VvJzVYYL6+gabqvZf6aC7j0sx2c6F+7d
4GxXAFy4M7QzEhxoa4umFSnwsuoN0FSW5Q0KbJudS7F6xNM8ulFmFRQ8OKdZB9h2+R7rr2t0HhQf
ait9Ekvxzhzx6JDo/pPXrLh9LijJ7zuOgmuV+uaFbi2f63lNwGYpxBYMCH313qNjN9bNEBDl5EOF
sXjEMnKOCs5grQH89UYgvrO/CN+gFdzbt6qcPInSl0wwDEAp1hBL83TuwYs+f7XYtFKe69nJSG36
o/+z+5Mu12JtLDyYsEU+2bQF69Qw12I8aQmWzZFA1fJ5hhiWsn45xfs66mfKzYfnqt124Qp8xoE8
NZUzi3ib9UU/Mp8WJqMkI2TQZevUbCwwzoBLoVwg87Itqiuj71+CuDOYDQ13f8Jw0c/jdEVuvHfX
4Dd6b28GLVXDFAzlrTk61qrQ9/JIsI2uzR3hmqPm6neHOgzbbLQTj6FWfJAo6QFvR6CGP5gCPScg
qIMlvmIxwCURVWMQyUaLmtau4iYI5349FWKXPQjUBo6Hq5RPnZ9cCA2vNcN69SwweW5vIXAn4gH0
eamYPgmLxv1e2kN7IMn9NDiI4GdMDxi/f2Wp5hKVvrUK6mqqkk65o7f1cDZGFKjL5vJxWA3rUC9U
69HVWHdHb5VBknmPSKHng8oSQkkki45AubgBsHNzjYbBsH8rAvMyiFU/x1QBKziNb32PriJXqSSK
aesq6D1q1FCdWIFl83Aw+TjiRQHQHPxwseG6tFFxz0MvajJmq1QTiJyo9zFhG9m4sqG71aVOAhoa
tngq42fpmpFDorfxfRtx0E025P5EYqAM3R0fHVslGoyJRLEfyHIumY1mCGgujAJw9KU0rySsjxH4
OBntiiQ7ioHw8iSWR3QFH+LNXEmKI1N95mhYj4+pUU03Gz45337PaPnm/r+XxKkCalDpnS7U1HmF
M4AqihGpHKOhFgBjcfrq8jhUGoy7skYuZ/lI1zTixjRa9jjURJ/1ZgjR7TFcH/QZjmQPnzpYbuXk
glrJWnj4cqMCeaTN44xRPEENbmNOonYkrU/vHb28r1N5U+hLYHBVzkaw/lk/amdnTDutNl3dfym9
TndL0kXvT0xUu7cPP9fewcr4aGWSV7+GdWT9Doi11vpE+IIHr+llPPmnguwGLmHQJYkfVFTE/Svm
LbShP+EW9LHwZgZTlRNYQXp5clq8LQq3blRJg5vW0Bu6rgbMp0SjynMB70vif65x+K6ueQCvT6JP
G93tLRGaQANiS2W7gkilo4Q9kupx2IxL+I6nALXODomwZmGwMbz/c6EYbKL7fZ/wG2L26yV3kti+
x9M3Sj8LcVP3g8E9VoeFbjrip8En6cjdIcFZZkGrDmT5RsiuRDZPO3Ol+ViBk7SOAhAVY0sfTP8Q
tHixrNftkk6u7I4mKz1mhGAppn/ZitkJz+QeBVMHxlguduChXOjEsH7y5S04tftiGPXVNUllIvSF
dxINVamiSph9JV10cw8MWij7GLU0w/Mo6G6IHRaeJBzGyqiTQq6w+PYdKJ4q/HZtZupsTxfV6YFY
Z+fQfzELlurS747d4lHWiMf1t/DacQ1RBG2IJMpEP9BkO2TT7gQMhMi47a5/aoK9WBKIPBtdmWwr
pcE4SnADT2ZDdWBJ98D4kGZJrNM5CJkCV4px4sqte9bXavaRk1EZ6rkP+nGg5FcjGPfX95gMZDaC
uYdAaYvaK0xsGM37xx/DdNRiW7Rr+wezqfiYH+teFub3o+A0K8I+3qOrDEREYmzrZnXmah6yBkQJ
NjeZDLdW5Ur8kKpMwcCkBxXoVZUiO/KQIOzRhjTQWA/S8wsttoEQT7859bOih92N/cpgpWEq87xr
SFJJgrUQa1RUInj3SvdqcWbeUpU3AMsyuw+0trtaQwojrcUQ3MTAgKheXdpZUEmf+nZ9+qul9tvU
lemcyxEy+4DfNzMSFSsrbQ0jl3KdKk2J2RwRwFz5iVhTJ81IIbIH5bBJi0cNFx6XyQSh884QodUc
I3jIV0eV3UCZkhnjRgcDiktAU1BOTQbovxDvxilVWos0JCgMZeSK8oiCuzpwMNVNG/b06Jj0Toh6
VxTk+CN498HOjg3RFIhJ3Q+YWH94JjFoJAZG4c1ITCb35Vl/Lu62m7yjRokdlp8WutZaeFVbT/M4
QiE2Ry+gnPfgHkAqITZoebhRzA0shqX/NyVDahoEiYX8vQW+q17grKlHDbJRvPxj0GOqiVFNfkNL
PXGBso0TrVLC45ZXYUtz22Baw0l+Fvh/94W//oPNuMhHYd7h4d7vugwgAYRJc4eYXmapahHF/pqZ
NDLQ65FUFS6V4pv2SQ0Nu9Cf7eDNARcrmQrV/d0dT2gLVmGqS7gPRnxcHGQE1RK56dkA/jf1N5rU
LvR7HAyIiYonHGn729rD1MW2Ux/DMooZVEu/5M1PkubL7D4rr98fFKviGiazCGgWUp4bikGsTerL
3iDtC+CsFakiBfFY50a8nbo0viMiLEJIsD+JUuXRtg6kE0LfWgYxupPd0ip5elfMJ2xWouh/rPux
z3s5ld7DGrKsNSE0Tc5AS/DiyZ4sBPGezCRcOABVSor3jU3GtwwtKkuRQhxLPMu+QXkjy6aBhZb9
sWL9lVUYDVyZ4bN2SwgZPSCR6O4Yn3ME6SCgiCKfbLioqKpW/OrkLQCrwRNRmGjaLJaMMmcRNh9x
aDWNXIUBaLEDJ+Bi/FX/RVyOLCpk+clz9eaIN4wWI9irzO8pKEK9TZvvLkUaob6E0Zi4mK9jDIhO
gDH0mWiIXfUDqvZXUBj3E0EMd9Bff/aI7jm/Hfwnnb4UU15DfWln1JmRiG0eBa8+vUq6k0NALeJi
Czde1meegrs3JIbJ5ftvt2rRnQDc23oWILYRV02b5SMt2i3/toSRIRkYXjfE5XikBmEdI4BZXAmc
qDzl32GQWklR0Do1lkDBfHnLilKIyI9zes8J1CGF6V3lNiZBDPWx7ayk4VT9iYT8eMGiIHqC82x9
O7/tPjfrVC/0tNb0+9wkmDWoaHcGH9wfZOtW9RO9TlnTqWjRHwhxG+d/6zcr1tzbJUCh9ixw3m1o
Y4mncb+RwZTDc0N1I/YdfbXD/Ap+FjHXdTjTO5BGWtZUGVqpbEmOBGKx+NAQIZKjfG15njVzMvAh
ao7MJNEaEDyvpZnrGKPD3nZZFl7Rrvoh+CdPwb30EAf9qKrtsiZQz0FuQ5tpXYlkENsQrbclRcmL
c01gjW9UeGFVUAd48DuNajB7jh0d+Et+vVeoPMZOvJfVfPbYxSSPmVC7sDe8wN57pg7a5GJAwCdj
PRibxiYzwnyuzdVHeRULq0oRdLyDoiXwe6On+8N+czajaoBJ8K6g+Rxna+chw2qU6oNpvgmus807
pdB9x4CtJGdruEu5CLc4KzoLFyBYt4YIjRsOUo0nl5PoRyyyijGcP+9MvXhqAENNYQ7EqG/CRpW2
y07sjIkRLxV5elDf2xkB8hsMpjCLBMWNQx+UF8F0kyZvmw6ymQ8E8uaeRx0NV3CzcaucqLr98if1
E5opRMBaZZawXPLCX/1ZmCJuaupQCgBWxRBzNBFZc0xGcP+I4eCfgtqJkZxPBG1twVYuv7eg0i5c
cFpLuxflDEeZzVy6q0xhYootyuTr3GINvO1U7U7Cmawc6MQC/AYZOPo5B9iaf4HaeVEy+eyB9yTi
H2dzlKGM6Hchgysy1cOPmezKSbTdfeXaTSz689L4HXSL6R2ORJ9FcPW/Lxv4oJXqhhmKpjiGTwsu
Wss3xX4Gt35JOzLIH1mimaeZa02QlRK81k6pHjrBd4ch7T8WE+KrvrSr17wors+y2INp0FHy7fJo
MC4rj4fde4ElRAAiBLWxx7fNXEp5rKFPEIcmWljHKQpqxkjXgmOLbvhZi3Zbnu/fX1gFyi+JTlQn
vsKamcLTXh3vo5t8nBb16PJyzvBgUBO7LHqMCzn/FIOx6dSjkeM2uWvmbk31arET0nmyMwU5dkY9
SVVfPY7IVobJzLIpx5/aT+cuXFmskPx1N8ts0+3Alo/xnWUP5fzY27+ZgFrcDhBIYfwI8WiQHGEP
DwbokipaFJI6mx/CqUqNT1LPDk/2mHek0HrA0V/mrJVMwNgVVIhmHhMoyqTaUJ+WC2dPPDkFGOZZ
QVp4v6cYUt1FRHdWeDUUYMAVNWQol4dtnNW/ucqJjn1jjty97v2IM6pRGZiu9tnFrfSjCggeUEcb
4ZkziN/59tFyhxnoI/TKvmEXV8E3qVn03reIrvbvarhKofcR0GjLIAo4PdoCBUGv7YH8cHkkukDA
ak5rdZrHgLEh9SYj0L7A3kxre4/CEvUxNURB4LfODOpoTH9U0K/CCUKvkCIEIGm13kBKfldhnS/d
EyEuusUfadC3PWOCihVCrJVbbfqESZvhP+LCoEMKYeBWJdr4HJd1bIxPd6Yr+ATFXxSQDPKXcg4X
/OZwuU5rBn0T2Rbn/xloa55F/qzWV6CXjxz3xWBT+nUGRZaLKrqjgVmBf2CTAfhEecWiQamTTIYp
kTBs5P1pTS5k5dsujRAn8XKvJ3hurvuLWFUvUmCAZz2zSUiv7+lLkIPJoALkeRcJt8UeFGJqDT90
yywURW7l4kcNQl5GGqM2Im4BsEzNxjv9vptlG4SR1tIzFnZ6BKMtKPUKtp33ref0fbyBBP5wOdYl
QsJKq5n1MoyLQMRmX77XVJyaVGI66/WL2ftcAN5WwDagcMObGLCLrPKuPNOpJcNVT5zeScOuhF1X
Iha7L8NBlB4hM3Jt2+bxpbvkAxr/KDt4WZGps9zghOsjAmu59LopscRdPsw21iWwfuIvVw4LKnmJ
zpMPmurTfWpVBIlNMJqALw6oumG8sWHN2wIaFQsOjQCiV9K2Ex8mxcYXxxmwXGdw20Jq59306ER9
nG/uWX6YI9y8WP1JkL7oNHerfOM6Z9WVRkHBaLRULO0X7hzGy7xyJRN8ilzo7hBLWm8/DwoJPgWm
TekJnJFw6OjauHQTcjUQKJ5TJ/hWl0qbeKyS7kiHoAKiXgZplf8Ky/AbUP8rnH+rhR7QclXnug4i
XyIsqivRNU/8JvWZ9wxNJmoZ09fudDYVoC2jB51hL+ESenkPl4cUv7y3Q3ZSzJGdnCdp4eDfT3Hb
Z7s2z4Z4+5B3mdFZMFGHm3RMS1E9VeUq//PtaRSEpBsYRvQjJGUamwZfj9CRs1gZqUagGhJDzvuD
WXexCzNJ2ko/pZDURxfTAvEPgBtg1/e9pIBYmTPwNu89nqPaU60zE/ltfie1ieu2jON7mUFjKk2K
AFcLGRWaYvBemj9Q1VpZ0PVQIhQGrmAzbdSIp3sYc2+PmOWPMaAYgeVHl9CVq18g2pW3kBB+Jytt
iRHCeC+d4liIpmPbk8DwOO4QTCZBjU5Lx8gMxWSqN3Gt8m22qg28ObMeUU9JzSh35Mpq/5iab7bW
QpoI4rltLUlHoMObClpGQE3qqQIvjihw1UmzDDJbyLqeYqPZbMYRsyI4eGZ/e5McIvvZFDnacFW2
qvr8BbLQP9jzd1sFADR6J+InY6TXbW2m5WJ//oE14mEG+bE0upLP6R6jnD/TN+RtdPdkKDIgFQY2
o1pUIwDUJMhKUKHSUEWC03L7eEd69fpzt4zX0xq0e9NqyVt0kIiYJC1TVrf7n8BR6MDv0rJQtVEL
kKVQKJPZg368A5PjcBSvSGXKq4PDZm6oZm4F0lVQPfIqoItagv+2WhLHz8/Mc+P9DyPGSyMOpoC6
FyR2yBLBknuPZwIp5OeipIQ1uCYSWP4efHWJZpqgESDHnGDFduEi0hJGsLVzqmfy0wWe9ZZxqL6A
10VxLxsJXut8J8EFtdOVeGobxXDF29jyL4B/jsPBnj/+VyvT7yFrIZDF9tX5O+lWHj2/IYfyJ5V4
EhDYvr7tYsj0v1FthE76Bomaz+CKjgjB/B6z4kxga02VOc/5i38sDgu+p+zV/sJ6SjjQ34S/X9jQ
3yyJ074JxvyZmGgnIvAGtYeZSvTlJVPP9/ZEBRrrvSMEAIqitpBRzchu9PY537LeQ4aUewL0ASEw
SM8+9sGoxGbpOkFCGkbcnRdofeX/BX1zDZtJHIpAKuMo1EdFRqm9BLRMxU8V7s4pUfd3AEablyc4
jEYW73LEwCCdyZbVOz6Sgi5+Pl8Tk+y5LMmYKFRHhSAk7QWCkeFdZ8KzsI9/shLMBb6xBqjQYnS0
PfY3+Dg6+CV3LPbmVm5lKBe2CnRzrscaNt/3xU56+CoXW4KWIp8ZjtU5URAfk85B+LOa/0bAIXbz
4c3qD/L9xZVQ9i0Uy6MbAaPZwXdG+i0KU64464SisHcclETm31sIic1tLx2eBB3fMr93M1jwkalW
kVsnbpdpzI52JR78aWc1CQVPdyW7GZzaMVhNLnf3r8eHKDJVxcVMpKGgi6kitDekhk0vBcad5e+O
Ml215AkUDuK9Pdl+z8rQmDbo0XjNsAUAqZM5XvHjty7fJg8UhywhMgEl02tIDujddjnVxaEX4sYB
mnTXpoxueDkP+7QJOq2Q9AswalksLumPsH+s8mJNAsBLwlYNMADFmlxKp/vwElfcTROHj/P6yPqE
gr1Ze1LmjKH4rawCJ+MFX/SV1CF28AfoOSxnUsunFfXSxQcyrOORIexFNi5upkS01GHpB0XMOypp
0zUZ7q6tXjwr5YaqGbN2p2207ee1Bm1z0+RFQIF+Z+e/5roHKzE7UjMmDwjYgLt6S2A8yH1q7O3x
N/9+8EeeXRhwhVOqWm27CzSAaUDpaB+qfFdNUIqH7JRpsazg/Kvufo+ALaQWWc5xohr8ZWCwOOzx
1tbOIChUBlAV3oHq2oixCJ/hHvjl56+Y8AxSZNm/rA774K+T9ozSdRj4nA/xOxvGEjIYsU2pTSpB
8HNCuDWYaM2obKt+Qye/lfO5Alnci2OHbhNTy/P4jp133d5V4jzVl0j49p4UjcInV8Z3X+HNJ3kt
V4fnnLC85X+o8evRKUvXcWXTSPECTG01OhFabY2C0KATBqCwBDH/ZEHWFg603SD+FOsx6Ti0HYwG
DxcJwKCbu4BpkXR5E2VvwkhweAOY8njUnTkWBwxwDgfz6fsFu5aSuPOyeFq21qvmls0m1xH1CXBe
eeaYqF7Q8SF0On0oSrxZLAh07Yth3UgHFbbGTdYHaLXiD27cfDe3eUHEk1FQcu5+jZ+dCUV2f+S8
pesZhRBwLAq4i3nOagm5yKaF7gQWXMHmwgznKTzNyfgk2wt7ZVGk+BM6Hz6WKQsDm/du8ZPIGKFV
IRf072+be/8yUBTk9pzFU5rfgh5woTu3r3BssW9t3fYkZA/KKQyDiAy3EUPQAHraT6nyLOiIc3TM
5Ou4UmWw9/LauMtTNbg5grjlW6RgXH6Ogg8NRSjbFMX+d1LOTLKsZ7Ug5M65Ker4UUNxpE9yu8nU
tLe60DfIMJIbgmIo4oWadVzJ/PAKwcTPTqMiyvoypNM77r1Beaycewo/WG4kjacpFIyHQITeqdea
777eBefeuE6dM6asldeimbHVkfv9mVRHDXRmhXK02i1vmUoQZwmSeMJcft8WMzBBQSL7fT9sG7ef
frhRis1afBvasPhc/BYKveR9pnzTl5BgO4t+X1pJzBZE+N+uhSaBw+g78MysZlAhOGopBn5lf0Au
dqKJoVnvRrAPfR4+H6lAJYtQYjma2rBGHIf2KBtz9Ln2OvOj6vq7EeJq+38RGmpUU7b1j30QbQsa
GQlwFozoJsi0Q0OziPgAJWJP8fX4UZPRlpqHSRd5nZ/MpJezUbC0LkDuMoveeRibMOVakdthXgNP
i8bTtaZIcmykVlnjb/CBlEc6Kmjn5yjS3DcT6aXBf5NwzwFhWlLFhh5xhSWqubFcnn7CpVVtlNAc
mzIWfoBkF44xY7KRACblaC0Xbqf1HGyeFK+YqfzW0mk06UZEQLeu0blRi0gayZ+YUh82NiSODICU
MXLXSrujProT3MlbjBg+K1IWTzPUlhaxcK21IBkFtm6gTCZv6PDTRsG+5GAx0s8y+X7gwWd6tQgo
1f3fw5qrJyQn97Rp0pahRHw3hBN3fnF/ZnWdsytBFzhNxHtxr+vhtHHSwcwBwZNydaRPyKE/rSqo
svhTfGBQBP3In66tbuW2UQuBkTPDiC/qqyhOGzm9DtYLBWQgehQfyPi1O+hi0D5Ze5IA/jVk6UxY
eGzevKflQJHB4TJ+QYhM+aRLf3ejTDWKQXh3/dHlpJwfS3h/TldDebt/WnBSBFiAoOr+M9JujIal
lbJ0WXP+V/P8RQtibNNc0Xy9lauWjOaY2Rwn70NfmKe5bQTHPnitHwIF4TRMb5SWOo465QSaSL8k
aNTOZWPUDKTn6OEzNwBSzjCEC5p1mEkR9RskPfOtxAC/UFtTaRgrJw+tFJ0CAudZ0gl354ss6iH7
vPaSS3vdrSHVVr2kvDm1IaQ50W6dZFwfPNhFbtp8wLoi34iqrpCLe67d2fpMmY8d/NuoD4oOYkPY
QhdiuER3uZXEbUFz0r+bYDW83HTAa853hcF+BTdVC8YI17iDIVNu7fM++1lGf8WCPHN+EB4Kowak
1JL23RJutQzvm/3WPn6pGv7+zoLwK/RRmQbFMUWq5UhfMntnzU6ropLigHPIXPXEGfqr98OgCK7b
Wdl0516tOxH/TTWhJi+/zNAX2y21pJlkFb3OQkr5TT/f34JpEgm9HxZoUVEfOk+76Ugh3aWhDVVi
p4B0681RsO/ohSOUq5A/w05OlnHgHv3N4iIHjtz6wwcQu8idkMwpNrB0wbxyajoygZZ3aDvOmU9I
4HBc/ajGHme1zQbnZ1ZE/G0A+teJcbaaAY/YbzlKHpGNokBkw2FsKTHn/QBSedfgfMqYtvAr+W5Y
luVIf7WL79CFnO6+fNVdNlVHnFPfyJArC29DwoGvw5NkhOqPCQuGuGGRTYPsltkYXd8MoMjPhwJo
wYvfTQ6oaBzIPfOttEkQWXaiUuqq6Ej9YpUqqCXZvjuh1hBzHDHv8pVGilAjw0hz0o/GA2tP+X73
acKAZVWXAR942YyqOkIzyVR1xZBievuWwPUlC/X3+kr9J0+oQn5fSpcKm/nzZ6S+RKH4lrS1vNg7
Vlf36bw9Pp5pZOzup8rutqjahkfgBjOVKlx02MZ9e3cDqJtL5auIiJwNc/qj9En8xUjgfqrr+qq2
Odyi6L4l/GJkFKvE0NDDO3Iza36vBd1rqJ+mmjBPtzojiNUbVmB6vedoP3r3tyVwK3x1DvMmk+N7
4ALLi0P5Qtl2GDErmCdCinQ1j2YJ1peCWycZeudI/CPlAivnFy4UDqFXkkHjqper7mXFLKKZUjAi
py+iozW9Ik7P6uuDe2XWU/5rVyQ0arb6cyBgcUs0/HVctDlRFxD1AVy9Wo7xUujMGnaAq0eioW5g
3zHKG7nuxfL7VhIoS6B3EF+F0ffiZnvaKOmi2rCKo2EWDRqxnW2sLkt29RI5emVMM3DNn6lzlHvZ
ER0Vup6pfp8DieHDMrDnCTz0kS3ay2oi7Kvit0HBx/qpVTMyoHsN2LiaBiK+b1XYJfqAv7LbQ53f
I/o/5g3bJFclyiDG5HSTKfe8nCXfiqWnTX09qIXVhW+4lng9mCdvTHeFnRBUszpWRjnzvu9UF4f6
PH75GEx8Qm4usLYOAB8b/kluAlnmoYz6p4PUmTb8z0cWyTEkA+stiiML+yMcH2vvZVEHYNynqw00
wM5/u2BnBubFLS6TkQ1CG10T/qAM1NoLHrFE5OpJMTOkv9I95c92WpYCliaTiILKKyrL74cKujjg
eX1vDUR2DLONCpdncw2bXn8gk+yXnsWfkbRobssfXywcyPq7JiDUTjt6NqkQE/LUjcsXadRpo22b
T7so9rni6VDaS8Om4x6xByO7sndzjAykqMNuR5jbYa2mYEKQ9X5uGHCirC6huXQ+RJH4rtI/8Bsb
tFUlQoLhjMdqUtZGC/B7Rb21lkimITyl+FYNg2gaxwbAN5q/3A+sZS2SnrYBxOtzpV6B6GusOKac
98xmGqwc2jikuSJOyhJmzLU8+TiNYJddO6rTN2UqVxbiiVmPGw1nOC4rrpWdx3ObECgUZExzLvDy
0RPrrbDCG4pXBy/Y7sYl5kHOg4dzGU2szZqfzeo2Hvi9fh225cDgOY/p8pIaawdlGXVhq+z3lAyk
seULVbl9SWAqkAOey4zw10/ZD9JSTJcCwxFQ4Zi+lXykn1NOrs08S/KmCGiWwrJlEf2lLPy/jAQm
7S5OrIRQTppH/5RZcwdI2YDV8mjJTKwQCCRKtIUQccEbRQnj0byOW1fnI7cJUkKqxHA7GNwEt0xo
dxg6CdZFSUenZjGvgOMmklTEUk37YTs5oFxryyETrKLmr36j29Pq07QbqwnRijQGUyMlr+ksNwud
ItvhU+DTtc40DBt9fmdyOhV/LCB1cXagNeiVSmk/KzGdDzKtX7QydYO8/OfjM2Ic4U2nCeQT2DFG
pzIBtUwhDv4+GibNSWA/lVAw5zeVG3svpPJqzlmp8u/pZzvzzKAKu1qqRDb1ny8CxxBSh15Nb3cE
o6Pxh7dvoGEpekhoSlFjwakWBf9NB+8+rgdD2/CfZSGi7Lz7AI4jsRHqTUwg657sve19bvIQ4EAK
JuViVc6qh/3AmAjp5XxqWvPhsiZb5nnFCong/1LTyGHgdMr8lMukXudTh+r/rt+gv7cPo5Mysz4V
oBrhDx3110EiZBeMq3As9fLUV/yM78TMKHvE6zB/rDiqTWNzLnccTftkRX/XYknZQrLeUmF551sr
n7/aX583zhM5+VJd0ckrloPYk0gPjuCllO29Pf0NRjj73LwVcIedPgT4sJ1Ho/3AyQU4Rq1N8E9t
hou3Iqc2lzEek/WVpRYQAJcTQrE6J3rIl1NFsV6iM5TrJSqaVNRzhm3wEXOdvRi38N+LHG4q0kvQ
lrVsdWPaOQE3WjyozOBkX5VQ+eUrhzvp1bdwFrR0rZnX4e0ByvkeAQSA7WHqSsCL/DbeMfSqnLeM
+FZTHZ3yoGDIs9vezWbQ29Sb00uPk75efgSvdAv3BK62zaC2IiZlBbL953xvp4jPkMtnni/K4hjv
ozjhV8DMu8uRIR8IpMCSpCJigoCzQcWlDq4XBKjKYb0CZqwO7Q7RRpCkIPA4iN2lMFm87/F+SJl8
Hd8uygDqeiy2FG3IZSRgEl8/LVAY+PlFsYw9TgE/6wOhXS73a4Hfg5dB9sw7B+yEvL2Rzg3OlJzD
MRuXs0xbzzIXgY3VQp+Mlj2QNGRs4C83hjWRyRQCAlX5zJCF4EJGM5Me3252z5502OuV/p+u+18W
4kxkhh/rmL4cuQ8WHGaV/zb1rXuK4A6XR2ZBs7vtMuqtbKzMB8N5UuYlHEMK8EUQCRv1UoTzWrwo
GjUCzydE3L+dy/4lE36vgsTRMvrURK1/RKkz0aNYRfIWdsMjoROAsz0TlOKMnYSkAYxGX2MK1vIv
GgS0Do5drizxyi0MFuhCMPvq+CvDQ1yY4NHECmfjpOlHNVsLw/+N0iRUZduTKimB3hKfgSWTZQQ1
kY0HVvhaaBbrAOsfJ5VM2CeCVUfXCl9Tk2nqlHaIdSvt9Y1lMA2gD3dkhOCbRvnYO5Gz2RgbsEAH
F6TOCz7+Q63X6o2OMqMugGpY6qnyqmioc5IbyjReAL+2GGnNNvcDO74KY2Hx+TSU4AHhhcEUBHl3
vBclGABEAf+zYL+ZgYFflQqVxV4NmPZWAsXtLJJQeuPnQS3EummRtURnQidArjAjAlT03JgnYAAh
l03ZBWtqobRuuKNsSqDfkL3/rufVUzagd1wO2/In3ZCC8DVEbf4dM5bOJ8e1RT3BwcwykdAUBRfN
DSYvW9kgIXa4OmyrY8GaI8ZrYGSL7NbKCwSq7kyhkzVNTHqjls8Ib7/2yYfs/ZN4nEnfagXj2ZGs
o094g0MqbWd/LrYcQwHfQiNNa9BA1mE8Q3nlyX/DxFw/ev1OFtyiWCRlfgcpDyhSfdXLrC/ym7Mo
sdkPOcbUOei8UGHv80zoBiJk8SYUPnjRXxEPbDh+fPQABoRJyNsbHDhJEWFVowfB7tmA9iRHY+ij
sam+HWMKT5ZesbQP7ZPFYzfMgwUDRY4lbwADQMtA2bglmZz5psEe9hXZFGVzne4TcdGx/IWOzZbc
FUVtazhGIqH7+hJkcSiJF8ohy5BKW+Oinbh/xCUHcbop8B6L9HinjPp7ea4deODJcdTjQTyKi7gQ
L0lkvD86cC8GDKwVWvM8lMOVZEHYqr0tbEKyl+gZ7IizzEYZLDzwHsoN1e9L3h5Rq4wHKOoVIgVh
fsehbZOZt+6VhbZZiwKRlY2g3zkgr5ohNyPHXqfygthOQ0KrGpK1wNnMVPx/eOz8p8JkelvbL7cP
E31YdgMme5PfuJJdXFqaNCxasa0AqqbGHC7LCLzQOiHjInWCwu/nzRMzI4eNVxFfSwSv6Qsc0WcS
od46D3wT2fsD15WivAX8ld3IrvRaUBOSsgKKuczwM+xjlRrnIlmGaPgB+92eL9ueIv9BP2JowJAr
zg/pOdDoZftnnE55826+nc8XuA5UWhdET/IXyS/nxX2PaCYV8S+MX6YgxtvrWytl/AXQ8DYBgybQ
mNRiK4ofNfce1XF+qqaqieKRE5dPfhiRtWaA/tmqyYrjo1OnZ1pubZBJs45YFtiQQyxf5/7/4DGe
L6Q0guxi/w27nSQfBM/DwTexTyEJKaXFo0Jq5sZwtuqf/xWkWzAdhPR62K+fkrS22M5DA41CQazI
sEStnaviup4TqI/YcGgtdH4DrKoNST6f1DSPIB0kH/1LPJAyN/Yvy1MDDLdzMTI34jYlDtSPcuxe
RYBd5a69O7TjGCjg2dRCOPMwJIqB+dk24jv3lgVIBTwSBKRSIXqbRkm2e2IkWKsxx8KGEmdF6S2O
M6HcCHFui90LvzDS1UcUWsuzrceyyn2oXnBu0ozdTt94nEHV1HdZYjlaB+6bTg5x+UIM0bb/lbz4
uKEDlvD2BlGimy3JoDOY6/V6JiCsBdqXhuMmQIelLcbduQzN0+H/CzEWBWeX2PqyxeDHfe2yYd5G
wRfIp/YpN1NSl0+2wyGKu8WUUdFvArgf9XUPaio076014uu2SmUuPiF1pGod9LSC0GRXEYPzBpT3
ee8hvhldn3lAI7rXzpl9g+hSsEN81LqbhIlnhmbediRxwd9A+j0+pFAIWgIPFeDRkH4AysplQa5v
8Y/j2rkYdosVMzhOcKujrn0uc+tTMNPskLC5f2akMFHvsVIO5NVTghwczwX6uJu2xLpfAypGS/fF
9Cmckts+QiWNatdIVgB1d9P7X4LUksliojYG3OKIYP3WjBqIYvwKpZ95vRJu2ONMLMLhi3Nm4QHC
kQMMAQ8nk+BOdcFm/k1w4ZAvH/C/rQusOhF/9qNW0kmbzGDn6i1ssPUDos5E9s4P++szZckjmbu3
Wsibbtov30tba5u5n/Gkn7/1ylg5e3nA2ayBZS3CAfgxxMfqAlBqeRhj++GnCgjNxe8VUMjV55sz
Wiend0Br+mgQ+INwdA586n9tUjes5uihtlNXTh1sXTZ8Qr5X0qyxGMIeK5dGEwSRLcr1AH+vBAR0
65Ng+qUMmaHEPKbk+Mw2c9h/GpdZY+X+QC/kVbks+UPdG7Su5CqVMfkaC/QFzQTtiuzBdzEMxV4W
5vQB2wOIhfYrNBe4vq5nllZHBCk7PJB2VgY=
`protect end_protected
