`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FJ4SZEKBok+ps0SRODYOfivgvNA2V4Nm4x3TmFpBULJNDkazjb7SqGYbjoJTRzdNn3BJMSIbTPLV
beQgNusQMQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VfMXQu5ICoEKcIGkjk94u9u8Fs2EpfbVKmHn9BB/27Mx3CAovJNi2fFMe02mF8LasM0e1Zmo3adr
uKKydUKP3Af1hI30xRte7medPcTo/53d4J1yPrM8mVgtnPLjwpqbiwwcofjHzG+iecwPlbuuEAB+
iGBFjlddR3XwljlX044=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o3d5RKkkcch2rryCQntNN47+m2qzmNHjG9NjTcn7Yy/cCDnTIfblfZTvW6i790N6mU0JjpldRstf
+IKewivl5HxZdVEX+QrY7yrsr2Ez8+gNzct5A9jMGQYWnYQXovJy0nbJpEk/PPUWSC/uHoUs+njZ
N1H/SD4dvlbXertgl+mmKvSA9WlX3FNDXLR7qADgI4Y8JfKapYTvMHCGTLhEkLrLRtgPTnF7Q9+w
WYhHHeEPHoTGcUwz5pvJaxWzquqJDLibUxIp8/Wrne9zOB2zunsoN2tqP0Y4YjHpZW6YetZRtpWJ
k3I6m/BTuerg9j9KpRffrZDL+u2wyggbEOLV2A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X/7aJHQ1JQvkQ238iLFbwggtwwtVSLSxX4s7Jrnbe3uUcGo59bn822Pfvi66dRHyza/J7crYHRKR
4A6PhvSzi/4+4T2PHs6XCkQwNoziee505CfRl8fTD7ei4bs8WHPErRdp6t/6fPVaBDCIhRhJOKB2
NqseCPJm7a3Aonfz3zw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gu+w0vXmbJNmzEL17DxAh4yPrGjZFtv+dMTGZL52KOWBNFh5sPn4SDI1No7Q8gIwBySjYIBGu+GE
oNvJ/2c0/93PQG63etVxSBqWxioGLJ8NgjN00qbxl9mUlmQl37/XKukilcq18fFWYr8pVEbmf5I+
FmGYJ0zWSIZ+RZCIl9bxu+TkDOd1qxGxKiU122Sl8v/BJwOqw1u+4VDeX/lWvwrPm0VwHV1Box6/
yEl55GWoECECDlpKsH1pho1S6W7rDUneP3pNkTc/IzO0ULZIhyiB9F+9TtKHIDLdnkIjJfrmMT2W
ayU5iFnvG629eLxjpqg5LIBQT0d5fL2MU7N+CQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6784)
`protect data_block
LrWlzZFiGz1y8f7d5GyQVQCg4qlRnWBdHWmk4hjq0pjSbsa5PfaATAPGuP8jq7k9NHktW24WrTQv
2/zOxZyphO9mwtPAeWSdr4yxY++FcQmHEoh6qH5n4+11NGVrpqWPf9V+ozviX/w6rCKYS3AG3g1W
ByZh+3+/7BroJKRyTKtcdlb5o5MDoFsSY2jmYUJVHOBY2SnGfhHP64A1149H2uLIk3rgMJ1EHcIE
5lJUcrWk9amBjCR2g9IDQIqgOb3YZgtPBJmkBZkGb/QyZQLX+hde2ISiiNCiEwlDfzP9DZ1ta9Zi
Dj8GUlc9qxogDrwCTNV9ig29ZEqOYoElIPuIUZ1O/Lb8do3oCSZspqni155gdOV4bhR4sPjPjO89
FeqM/5c0tpIU4HBFNIW7z/SS9Z/x7b7vUYplnScefvCo5GBex8ns+FlWTwtV+cCTtn1eraJvtFhl
hYArPcIhmQurjcWcDJJMLnnDxedH3Sieiur4e7mw4GcDRNOxH2Yg8QrRfTkX5HEIMf7O0GSEHMBv
QHDOBPvE8/W3Kqu1achunB6LNPucF+pn4qCmZfIwZx/t0fBNLAEO/ddMknYEaitsSpYR6DnQzV/E
K6es3kuPWkh0fSZPtO0RwU6mM2QwcAyn5vWO1YTpW+Xr0vz2TH5xMR6YdxcWavqiQgXR9afeG7Va
StcUy6+IyBDVlvUo2sdoQsxrf7ktyd7A23JDY2klQ936dZ7lJRYWTQhlcCQ+hSBfbBvo8g8vXFAR
Z1esw+iMsL4HeMBrQiLDpweJsmXwZZD7L70xVe1GhEMryDXpLDNfKm6zR0HpDmAFESCt53+w748f
3dMzzQQxjVrBBmxRdFkgTnVFAYsKoDHnlILPHPNLUklFQEoDQPR3pizi5laPRZbFCtCKrFGud8Xo
QGCaarvhA3H+b/vPl9WA9cC98Jk0353CjSuW2/5dwolUlvsmQClPCm5QWtimvDjJdaN3+oubykPq
DHDy4yHm9gtARFIICeHisLxzfUayJR/bv3f3+XXRKXNJzQixfyasyeBaG0OJmB2Oa9kbwnNJjgfA
WlppOGiaxwDOqN7XWZvGoOoKNfucQvHWzvQFc+bd7DPwzNnfLz4H67RYd9gm/elZXDtiWvOfNioW
0hsKcSe84x+T/CWoRlsLToQ6Dq0ArNX/HSnVBe6C9DCMGF3/XtvnE8sf16ph16AaoMm83eVfN/qL
75/DWhev/rOTWtrZpZPS4on1k71V4j/CJgTWr0/OfYE0stn5p4sYWIqLkFZ0G6xduyWT9uQMkPSf
Biaet0tYYyTxTiNKhhdhTgOQqO16goF6NQlybL1/FqejQag0AwW9nt/VEB/MhqWY3MwArWzfz85V
rtlGXnMiI4rd7xVfAgItrDoX1Db93APajC6Eh95iMPlKZbXZUpL7mhDUswI7I6vNWs/ExB1rFx1J
+5RQIG3BXicidwPBqpOeUD6tMuKDBfgCYXGfzHMBV3pD28guVrGmxchTVd/+KQMKjI+O2pMOOnhA
ryfMCg9DiUspleKVnL4QK8aXqBzXJuGajT6q+Bx20w4zESWOlH9vsYQXNBgit4rTDeleyQaCS5hw
vHigu7hJ/9C2bChfDDdD3ZK2I3hhw+ldzEMXB5XX1jjBuH6IBaaFbQyp5NyPCxgoLyUo+5Zi3oB8
vNCqZCw7qK564qgPK97/cSm+0lpJW91AdUessTICDR8qJ7qR5xvX30jZf1ZBEDRiGy32BWT1k9RI
UFFe4Y4F0x5L1pmlUOPVeXhdHaZFULA76M+nYw8yPtsafRSvHbmF8B+tEGOyO43TPG3Bmpu3MlTF
K/xyvgt4r79fmPRKSwGFCx9EBux+QBrAzKwYGlGz8qVVUsh0Mv8lCZpSx+NfFJyIpy1OQPPJUA33
Lh2KU22KxBDOteGIFAvafK2fJx+E68dqXrB/5Gx8r9pkg6SPDZBbzpkHwokmnT4Z7ArA4eMS6l4P
tXuaSORKKwCIJqCmF2cDOY49HJPItRnYjX7D6XE/ITTjq2iwVIWK1OC5oOn8PLfQXJk8kkN9up4R
F3iuMwoNsicgruxxoEwx93x2FSQo55YuMzj2cD/H/ujLjlLzl/BYr0fneWuxLv4ptz+pWryo0tpw
/y8UYhrJ3KeBCvZBc2WK9f54bqQhGTx/QTM/J2Mz8NP9w42ldQ0v3Dt/h3ZVdRpROosl/mEpIAm8
tyEQWZ+5VafrS4tVAA1iGBrRtSV3nFFEPmjBzIy/HRbADbLsYodSQFrZu7wmUt0ExK7kKLfXytR/
M5IA2wNuW1nQqhfN65HTfBBjig9KaJAyM/CaI/prdIYE174oW3SgrOAbVzWJgUiPWaL1d+ERwbVJ
rXmxuGf5SjkGRSGOlYQdYKpWQtYXA1wUHxGLCc2HAhpZlXYJfPCh51GSh6Vf9PiztL2DtAYzKqKR
T1drp2ngIbK5mGGJ3S+JOC5wXg4FT1gl9kawQeg9guT4qBaZbm5A/M9O23TDML1WGL8IZ0fz3XdM
Pq96CdpCXZJQLbUkkHMBhk/yC43YKi9P2d3hz3WBdPVG2lWKuVSXP16IrXXha7Vsjdhgjfy1yaRg
ZyBwctoMTSjUeAHKjaTSA+dPK+Cth3PDPv8dFnhgYxYxYQsCi86p5zT7WumfPXZ9IHz4K5aPWtYY
AlBSF30okxKc368f1JbcE1BLwf9WXWbKWgi7/4U58vNzRmX/rV1BBNZk6/Y0aTSGFFfJe2IYX18G
D5sZPf4U5biraXdIjgH2Ah27cLD2xeGlgUdB6Wu0XoKYOq3+Zswsg0MjWn+knkkMq4x4ZqmDqaC1
cUpM1Z9ZDBPzGRSiZXeTOlEOnITejI4R7/kdN79YoBy9gGFyIBRfbCg3af7IXq8hTc9lYYM+CMZ9
MVEP9676EMqyUz2gZ6QCe9kkKXrudxW6iQlOhg43qYRfDpDt/KvCkrNt0wzjuxvFBrdiJhKOmLth
1OdWrRGEyX/AWghiZv37HpvthPpaDId40VWCVtZLyEFO50tpoZ9GLjPN5HUKlsDyMGY9tR1QM7EJ
/PfioN35Ikm0vanM9kNrqqW/6fnkHB5kk6poU1x82ICmZazWF7pDqqrI6mrCyMnhn0C1UdL5ma+a
YjNXJthp2Og5/zhxr7saiCbixi/QqccFfcUsDgiQ7eAHo2vYeNUYxpomhWUGijlaU6XK1rdoDE2Z
vUz19bo99apjQq2W5n4/i8Q4DLGmdnlyDp0PDKsB0R9jRLP6KAZCwjJdBfBYiC210V/9jahhIKCL
SvNfsdiaFFx406Aq9rxFDRCWy6kz2CE8tHi/exPwnDD2dgFN+DL16xXfyRqwW6TOYhC9UhcrNczl
Bv8iWqKdyZh6lwmqLGAW6ZoMyM9ktRiv6LQViwUBwAUmEn4VrAdSbBuPAdJjXvpPmejtxWpPXrm+
bjx+b/SY7rDhe5gtejwE97ZSBMqBLPSGCsIeR0ZLyf0sOq4A32jINyUnLRDip9iatKXliyxkHx2f
wWjln6YGQiqFe/dWPEHX9WMKI8Owzs3Xt+DinWxtkaCiUxmKqNQfx9T6OKcAnRVHRqQr9UNIPjT6
1gHF/IXRL81CMPWMkhIfMjUG1cB4StfW+kknfHWqv4eg4EBIXbo8aWiIf0tZH0G6nyc1C85wUYHy
HDWcSOMNzPZY6BfYuOj1Mhfra7jyfJ/kcwv+qOW7JYzbGJSEl9X0i7C5d2G0Mk8QbFD/GF6yzW5d
FKO6XsptCTd5ZkGOjNDcO8mMOqIcxCLEi6zf8Gkwymqn9ORpNjR+98j9RA0dsYJSd6MB8Oq/gPh8
/T9O/dfut4B3o/T6LWlPIwUmHzUDe+geF3j6rqQajl6SGBr49eodqFsPoiTJ+by+1g2xwrxTHOLn
NlRmMyhe505tKwpRuD0rTnV7Y+0BFFA8N1Y3Zi1FrPnbPJKFBbAiosLAUhBPAYT++pmjymxfwPlE
HSpWEyYWUkptYJk415mIHd3goa5lpdqEWJpsr47lbInT3OAjqq6Uar6/nxE6TRm/7YOuo5fnysmn
TEse12a+uysuFR3gNE/qvTBrMHdPFxKo4+FiC4ZCJq0+kPHKwKVUm3YQfi0Ty5Swo1blAHPWLZYg
vwbFFWRbGzFHsvoqcM0JQQUz92NmO2DoAX7WouyUPZYmmGSOzAut+QDU7YgFL2bGH3ecX4kIUNri
2nuXW4oVfQ6zWaHMrBt39Fe7bnJEzc07QCCTlOONLbCnuQumXTvNu2Llwg7rYZxqrwFkYK8A+sVg
T8szpoCP2Gq0JMVVx3HnnvvzPtUNGElM4p0CptvwHBXPGUp0sX0+rmH86d/fomfb+w+bZwRLQuX/
MVFbfDGc3krXo0TiaPOvOSkz7VLSAxaYGJgWwQFknKWHKAL0CyHYeQ+P+m3w0jUJTvGNV5iV8XWB
NISnCLWZGMn/a+UJFEedQV5sDEWQh36V1mAnsf5LSCz5BT/Nr5bQahFRXgc5MAteMvs1XlpkJkQ/
TacW0ve70Qx11y/jVU6wg0aGu603bPoElHu/KUt4VaQaK3S1f5Le7eIgl9ahfwQaYZ9MIYKYKiLJ
iGlwxAZgWKwewWCoAK9+g5kHWGiGxyHQD4fFzLXKTs2B9ZlvPiWg5BED5FKHYvpNBtjoy2uRTZJ7
RIeKdRLvH+ruLQCCumL70KV5A9y06fNs4fr1Pe/AKH4T5MRJvAV5h4kj2TFzJFHV+RFT77zOEJ/8
AvF8UcIrO9QBRflgy6PYhqseHPnZKJR++fq9+2w21RlQXoXOuYlXsxJxYMQSYknqp6Zs9C8+H6di
YRX5b3a/FOu1KlXeu2ULQoc9LWe5+OxVXkOueElryOgu+/dZMGSckiR8MTG0Zxze1GG6pO8+iOyn
WDEU5hMNQB4TQT30cBw83AjwqKjrCYVOlXYpusNnJgbs6fmnAyXhye6+jj0ad09nYeO9D4tkxQfs
yfZ7oLgKhN9bwhglg1cwmYObg4G2Pi2/ffT6q/VGSLr1dqDft8dFAuwiEz/Jycf0AB4EARIYDc/u
zF8YVodazjuQTedvANWgzrHg/Q+6m9jslzsiFC9u01Yts4ItzKs0r3fU5tavpPomztXTsxNI/6kT
qNOoddUvAmgcI+FmtuUD+upI5/FKRFaVT/1EOKsCiGQmpsExamUu3dCf0Kul1brCdC6YodtcGvx2
sGNU6t3kh7E3SoIJlLbu76VCEOWko0sCD8pRrxrYnwIWP251l90NfRw7EsJQ3Tz6PHOlM+HJWxA7
Dj6xr+rw3kkA/Op6DWoEMaUBsHeYKJ5YqJky0TCN/ksh5gPseLcp+DRj4WuGQtChG6dRyaHYHm9o
nuLEebgLdup9KMFN7+XZMltkphYMJHZrqfVLfee3Q/qL48I8rKavMjmrL8JlbG2DP8v43vnUFzdi
KFYYJK7jQTrH4S5ZF9tZ1SQrD3niktE78ZQmrl4W0WLD2Evx1Dt8DVQObfZq1mrVn1Kaxg8P3Hoy
+LZiAAtIJ3IWMTZ7qzOKA+tUVjofLIjbALnAZAr8Pu8HhDE+lwWfG7xXJHvmOnEKjF9zSpagFWqE
TtTqYga8heUBlRs1U2XcRO8irQMK0x13kgUzDIc8mNYfB+9fO26fVhAuEPDm+m5XmWVB6eEd/nes
ROxkdMpZg/Jb9/lOChvNt4JOGqyYgZ0cGgjsVBxeyA+PV4dsjMv3WyA1hSly2szmCNFxr3G6v4td
meumTAzLmioPOUHMY/WF4dBzEbijQBAOeYK4YIBevhbvB8kmJJWy1RJqsEvvYdu0oU0SUZQKNXeG
vjtw8XmiFcUqJcLaTr7++HGa9OXrPVHeqW2K5aqRXJHtxnsyhoaZ+5bhNy/TX4VoKE+q7SsLL9xL
ef8/C7x87K97ljg+Bg1li7+ADXIL2Dqpk2XkwOLcj2N0U4vb5EHOdCzGUdjEJLp42NIGiwV7+bGJ
Gt/1uaa974KNgptplcbSO2TAJ+NjvGWpN7pGwTfAbJ1UqV0y0ds+odPR33ePcdCeedLVtbpSgN5D
tLmT9V3IKtYHaxnotaIzddzLL8Xv1i3EgcRkEOtCNhTfUzDGTT29UJpJ5G1sJKoZM4+w1HuY7ZGN
FFz2fgzKJpqAyFghXEnXuI53jDKVV/hGVHWTKg9rFmid/T1AZTRfAKrL6ZO+GNqASUr6P2WJZjBx
mXr2jfNBAkZgJFatgpzVsBhA9rQ9JquhtyM2WOdf61sIbSzmb1aPLLFhKmCbLbr9PHQ5yw5Dag27
wWw7+UES2oL3awVNAdkTeVebKMk5TGC8fb6G1av8o1Q02FI41/x9ihE+KSXsCfWxj7JkXgePjh2j
+8+ToHeFym7hVZ6BGpy1PZJpRkmohb5MxpD5/FWrd+2qpok+yMmWVuC4qXawqexTKqIry539zpHf
6/k+chxl/hvY3oOXqdiYiE6TiSDXtNUtnRm7lBUadG8D/sWpajeecXMwRk/+TYE6ytpAYwEHBDZz
gW7hlubS8P5vU9CiSkCyawImC8L7b6FH5bHLzg4pbD/6ZrcCpQrp7yEqEOYgmBCVUj8INlWnqguL
E5OC9D5mUHEGndYIC4tWyiY3kbxjHGi7oUcfPNY8PILKeOQll+kpfVWEZlhvO/eriImCO1GAPyGk
iYcgnpPDJ3+SJSnDlsBh1tAWO0G/uDYuJfSXTZT5O45CHZ+B4vr1K0m3N5fvCcxHg1M1/orU0zCC
fU94cLOBfffnC4VAeeXIXDsgB+qFZKrK/3yP58N+5oOLRFYTL+BM10MoeYyZBFGS1Mw7LUkfN7p8
BXSa/2xcyOKwlWfZo1RT4NLuVJhf5GzELso9l/X07Wtsx/2U3AZp+ZKYhHGmAYj+IWXLy6iDmDeb
l0gzeBAbkg494pcCfSYG9ZFe1c9caD+N0liUR2i+l45eihTTJfo3exLli9WJhFT+IrE4k2oDHTwd
2LEt3vr9aZgcW4avR+jQGzNnT23s6EXhhjADTjxX1Xf2Rvln86W9+m5Q2MGGZCPv7jWrSMuT16xh
jy0a1zyoOZJ++ZsTY5kslavvI+jYw9xzfxFpswCTkY6LJqqqh/RvyuBEulz286SWKevUAjHfmX4y
G5th+MS0s8vo/W6cqobWaEcvKNarECTkEvTz+NXTWaEM4ILL9NtqBg+7CxCPD7pmA/i1lkSNCZHR
NZahV2V1PDFYqyb3f+908ziz4vjxfu5ZwEQyMoKkV/iUBG3GCY273UjF5oU5msCE5C0XM3W2YmnQ
BPW9EVSOYRZHjVZ77dzEcPnR9SnTkd+tlxAXDy1CTHpJ1eSpHHuAOwXlrkH/zPPCXOOq6Bs5xXvF
8AgUWYJ5VoYBvoi9cYteSX78nLhgc3VnQNfTPnlJv5GlHaVubXVkH96JOCbbPBy7FtmPZUvkVtZJ
eszbptR+rkrLDBkipmjhnN2psaoQ/6TJMY7SKNg2RC4VMDcgqud5RchtJtrCNr/p3YKEy4tq1RF4
h+KMJRaOSxKX5kqLXMfBk5BAiYT4AqteXlZ8Go9Fub/ouwvsFCkUbLh1DmY+VWD9moqm50jmj0vN
K2M67MxEYcZq5rv2YrVjXLjYuW0OG7oZn/KuMMzgdrn/V4xrBr2KNt+JT4Xkc5RSNNY2jsCfyD5s
VvvBw5CY4UAGzvR35R9EVHu5Yo1coXZg7CrHou+2Y+zaBfcZHf6CbG8oTBwRQi36VP6nxM2ewjqY
X0wmT5dwDdeP/ITMkuFcKfSz9wTF7nvJvOinap51P6vdcgJTVdeGJHzOsdZOB7Zhha7N8R21PiK7
8dTeJFcqzdHlJDpXJnNkA99N7wc0W6XQG5dFhM08R18cFW8JfVtaqsTDdyfYYQzRHnsfShLRtPhs
ERyCbJOLhxqAJRSR3HvCocImKcixbUzQTEi5TaL6kDweuZqUFkQy2BfVohseVHM1DGWZ0D/9nVrI
zTZ6QH8RIqieMZUEMt4VIsqDoMbPkfWKtWg0cjZOZWQBMVMvrG6tn3K/oOHdZHOMGFDcuib3hBK+
4aeUGjNIipZhS/4YRnu4XvgbHuYWoj9EYqggdy8EhxveKQfGsFGdJwkZPDWDq8Dnl8gOwdZAe8jJ
whGXAVPLSXSnPQgxtil6BFNekX7wEEi7Y9gYlvrxJploanG5oa55pb+j5Nu5FPZWFMZDB9KJpF2b
3f7WHpDwUWDzX9nUb9b+sW231dDFARUIU+n7/UJl0ekYc0h0GFdg0W3mfwRxjQIgPbvMW58HAHuQ
7hh1UDZL1UG4Pdgj+NwOoR97qWcoCArnReI/uaKcrsBOHXZREsi/0IiyIaHlBcWMLshvTgMn0UUX
tTJUMm2AOFiA/LfaB1kRGzp1zsnbdYa2FsyAVxvWy9OpSTUGAUYjyruAgpqWMzTtQVsd92QJvBAw
eSXHlhTtKTrOVAPeSuj7TN7IItPjo1jiaB6+J2+5A0DrE/04Ix/rFQ2u8fPOrO4x6KmovJ5+w0ye
7zO/F/5jtFAln7a/tf5ZhkGvoAWYrfx1p7R4YlqlPbxQ9s81pyphLouh2UiNYdJx0ABILZAR72Fx
fH9LDQPNKAOtPq2pFRuXkqd+VdzDd85zRD+9qq3kwMHSW8QcbnL8ZRnMFGUaS7LVyjhelqRBAgQA
PJOebiY279pwC7p7ykFPf/vP2CA2hvePiDfbnIRPo6o7mWXjrdjSDI2bv4CR+i9V9sQrgrImruwh
ESPiMNsIKnmnF8RAiD/FxK1E8n12mN2lsMD06o21p+0r3QhEA9uJlh07RUdYSEha9nwF8pS/rlv4
d6iONICIFpuUD4Nfx4RKFvj9RfVm2woIzUtMRCkCZzYAhnA69UGHQXIskFGvR4zhcsMiFo/QPBbB
OJYjhs34vdHNsxL9dvZRjUrgccOnMGCOejgnlujqV/KBzk5X4WhxZ6YAdnnSnB4gJjbU4xTziQ1b
U9ADwXoNJg0qnyt22jH8wgazT1F8uYiSV+D0vwWQbkGn2CiSiozrOAvxxeUHnfpSidcgnInEELJt
lNBM+2AvmFrdWxMsjIASC7/TNfDdES3IlLf21aw3snjiDGjFh4VFJNv+T9369bwYdZZbEDFE22DF
FQ==
`protect end_protected
