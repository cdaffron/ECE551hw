`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NoQRsVX/O1PJ+Sg09cdnLT0eN8x/X0h7n1lxtGqvWQhCm/z7hdOdhN0O8hKGX+mOMK13PvLnJO/s
X+nybmKQ3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hGBSeQcrOeXAPGYE4GkGc+bG3KaiuIJ4tieYxzfQyLmLVt05wwMlgSvUO22IzJH/MjrLW+hyypqf
Lc+uNZbTQFJXA951OM/X0VdYLs8QL45AGT4+LHzsFjaE4h3jFV9Pc1kU5X586utzDtur8JiYVXOq
CbzTW9TfpjcszGC7fjc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M7WPOHol/ZzCAQKjv6IBSC6PoMqWzlO7s7zAoM15cUPd1zdPJ+tIO2SHOeCH9i0swiEGLparjZWx
Ivi4lApUiPjlfQo4Qpwr0DzUdTazk0ftdqvzfxWT98XkXSf5z3P+ycyDhC8k6AQEmBPHGQSGwR4I
HMblEITc1Wx/AKicp4U3E2U/pnO2RRY2WRh2XM1GE0bhAXX2QlkylK7/3xwK9VEH9PNfKd6aAq8t
+NfdyRFJSHq/Zf/RLcKe4LV9PkjcyXY8gZoX+6hVXFD/PIs2VvmQUk0m6rfuVotT2n0MVsMVI3xy
IR7ExSVaBwqPx6BT8Cu3a1grn9Pf12VMrG2raA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F5Nz9VN1GHSxpwBhCJvJ1cd80AOBhsQcwv77ccSGGbb6bN3NQmeBOLsu4CU9lmmOSHs+VDT+P0xc
+gbRtVkYudUBDAkFXH+u4kRXCubCMuA3iS6npgR58aKAXp5UAgRawTBt1yoT3Z/pAjwMhdy7pHhF
NQb7qPwL/cWhDD3NUPw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mt0B5fca008qUPt6eSR2Ksm9/KpUC9Tc+91GoLZhq4VVdUntomTL741TjVAZFpiNbZDX11uHLV1h
neWOYpA4E/cAIKNsU5cvBWaypvJUxEAER1WATJ0rk6QCXWSPjBx7Xd2vLV03R8PGkXliNsTCG0Tg
vZmIXqdnpJR66I8AJmqDpsN9sMUE1oc0eXHkrYbpweJrQ1lEPetLr5jqrVsQxnjxGoyx97Aw/Lm8
9RKDgnwMLEskzZc5cd1g2uFFLMTzu0U9nczq6HdeYCAIo7EcK1vALgw/H+/xYi0Zc/txCjt0G5t9
IUR04AExgziNCzPJPAdoNdnWZjfpNGQjM1+5XQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5856)
`protect data_block
dHCuU/SyYX3EmaXIw9DjGubWAqhYv4bD29Eg15Dk0mRKC2fNzlJdzfn7xYYTkhNSeUz2GAD38LQ+
5FV7/der/Ku1dFPJDbpTKhtwrHWOeOjHYKMp2JiHsq0u2Jgr7H6WQKOnHUiFm3kUR2cCpfbcBFGU
l08L/+QKVVz3CB9Aw+lOZ8hO79JTIDPl/zUEznr25+9OglX1uee35zWpldQwYY9KE3K0eSl801V/
OA9/jpbBjg2G45SP4JztdWekSReawpqOczjlpn3KjNjuS1872fkd3WD4nyHrBrKpZwlYOHnyXcwH
KQHqiZX2IeaHzWhlhmZUwccaAFKuLM5jLJJxx+SulJtPQIID6gA6mgkXJoZlLvggeRoqhTOo6TfO
VQO7MeqLH8WDhx/8w9L916fvIKm925ok85tjRmR1SOi+WXx4l4JDEQc9+28TCtH5LTd/iiMQLlfJ
7Pi23n6c2aZ31MI1GNwaty2NzvaJGDhlhvSQWG8XPOmyzv/dZ/JKoF+TSCZYbPHysef1BWKa20qU
02iWBgucl6fsnWMvT8iwZ/U7m7Vex0AyBWwlnx+l2VjfjhYoYrZgG0bk3QFoH1W03Z3cDJFWnh3c
DXuDCbV5DN5O7Cg5BQt+HFYbSpOqyOrLqHH9Ein7FvNH7bkVQPQWuYRW7SMmxgSZ3lL3ZESllu32
ejLKOKu/1lQaNzgzLbNu8zwZ+szlkIttvSb0xY4FMbuBHznCQfyHk0HDxJZ8UrNiTXUcpKfVGNGo
haOpQNuHTd493DOsQtIBJkN4uB4LVWHlTqcfvSGSlPWC2QL0mHo0H1oqV7LBZxVp1GiAPcdmRy68
g+UFrmt/nIoPNI9PNgOOmDPqUx6Xpf+mNuYXbFXkgEU89VzdROZrbakCVoVEVe3cFsANhfPsIm5F
zkNWkuMpwWc8ylbC2ORur0shnUcCvRMEtJ4ZG4JiEq6thDE0FvKg1xslYQNu0Ir7gENQ1A+6jUXl
7gQUBNHxgya1Wrf81xGQCZ6vD7a0I+yVZqapGpepyJWzckY+swtGM9tvQO2cEAStvbN4+tI/bq1g
6x5yRU/VeYs7u/k286MEo8AxRj9wlWUHi10uj9Q0kMWh61G+LWaxm8pC6igO6WjiYlyjmf8MF95H
GkvQg60kKdV/zGeVlZFRsv/1/5DwgttlpEUylMh/ZVNXEcgq00t5sBCxJ/agoazfdujfTy6U7pUY
fm8gD4RkrY4uzwr9xWTNtlDc4fRbJcnWWnfMeQOxdS2OPVUtH7T/IrxxEJCv/+flGsBRlWZvEYkP
slSkkS0PhxeIiE9mK2X0gxmOZlrFV5pABrUlorLk6QMTvfrRJv2WRQVaSrY22KG9oPQM05HvfeDL
7xvoqvJ7blUoiJiOveG5dNPjlItTaChvW4FxEDbMgeYcQoxpHo6jasgZadKw9GQxHfX8sR5svpdZ
PpvjUdYoGi6/wkj3KhpVkKYE6DmwmMTwmusKyz/Knu5cOjxOOLl8x43i1pnOtXOT95fq+Adxa0eJ
PFRberZQTVikNkCU0ivW/Gq4WMAOHdApUpDJUpRZ3FuQbeIa5kwnyCvr2i0GY0w3fWkm/pu/qgi/
i/ihQYXhi8NIz84cyOZhY3n9Yrfsffg5HILQhgyLX7H0Y6p2QPmJJg3nFEsrvKXnMHIRisw12IY5
RH1YSjce8U1YNBDH2OoafF3p1GMBxPJwPRIsDfvrz2g+36MRXg55fJ9gi497GcBpFPDJ6cqyNzZ9
5RtrimBfCF5bbslTNv600/LQ7BAq9o6a4u/ygvTUX1zpdqpYnIbGaEPh6PMYp+fsoWKqVbdRyeRo
NRZBx4NkNv7EzAJyqM6V0OnVyYnIHFEaw8hc9/TXJu8pL2Gl27cTKkhMCGBWxYsJcMTyHW0evzjZ
I4rCBzFkoY8gEmMiCKEFRoORJnCv1vnNiZDn2lHcwul3ktzLRr3reN663weJGgewrLsV3GjQbEgY
S4ehcTfcY3GVorcufWeqGdQ6EM2dpXYRWqI3hC4A0JlWGIyIh/KErPaja9CG0PIwQ+/s6oQOOFDU
kV1mnCM2NvC9P5NHg3DYr3K4ua4GNJlGVb3lJ1OkoaplGD9YRAGsOcPq3u8M6R8o2KuMrmAPwadI
GeDn2JDuAi1RqK/Iwir8Sa8InRLmjHG9w+PsPymlMlif7BNcGgWH0cwc7X99JAXKkWh0BPz+ujTr
p0e7Xiu0AxLlFg3B9xRqpHYGKRZMgfvDjvFHNpjpwP4RuULBZzLkqDpjxa0rDtdWzYrmAZm8KRhh
PKIwRsiHhdWRYse9ukyz4/p4X4PV/r28x2iMPzDTeaYyLU8dR+O3pjkdRCOlBEv7khxxqwscj3S9
VAtXyGvKYtTXyaq1J26dQwLwIUFA1L1eVFbuaQcXJNqsifA8QhKIP1pB//9P0sXQWWJmrU+22Ezm
3AvC3eTRtyhax8gaU1W4BN+U5AfVTnA1QyTLfEO0v+bY/RW1b9efBnc0oI+aFJpNK2LaWicpNamY
n6G+k9sKs/+UG6X5qW5k9rRACblmiFJdgnTpgkYE1fnTCDFWvdUkTQKQYAKbfZWSr1+KrfNxzWYY
yHBX4ae3qcE80toqIkK2QP2RzD0KKexCdZk5sHTfQ7WWZEM7TX3aEUMsPRV/OalS1BHtVw8wHeJ7
73iqjRVul2ybJ07AfUYFNaJxIX1HLFpF5XSLMEAGTkPewc5nqpDeS0XM5DrI72ORmDkL1b5+C6Gz
d8Imra+Qtql+Gih6e85oOkRwWWr6k0MVP9Y5E1n07wBr3nuIj/bOGTGi6s/zPKNoRG2cMtc0ODL8
MsGZfojyxGkRc4lOALO532yjvemEfv8izDkFKzjnqA7V+k3WnofXybB2Fpg2P8uD5cGmT5B+UC7O
i+FkbuNOMNQOJSWqOfyA5k+aq4Q+JEb4wb4FEl/39DfjyvkxAuPEjzRv7az7RFC10CQj2vmBDctU
X16Rm+WzuiusEnIXuPE4OVw0Uxxu9yn77bYZj36+rJdC5QtEqqxr7PLHvDwRS+/NvQNR5SVZwEH4
0cfh1NLSVFDlCV7QsypW90j6RoQ3ZCsTqpgspvvwi9ow8mt8LNSU159qTRjEG83Glm8hlG9MyMMQ
m/Hr3rTgwqytoF4u1yWZzYbeURDaKILSmDddkPTXoC389cd2nLz8pPL+PxWVi0XtxHGWdM4JfK0Z
2NYO7H481kfqy48Y8C4XDIfy60OffXH0Ukx+U0CVrsxUdeqvkqY3os29qXqwkwdCbQ6caPXxxd+b
N4B2I0R+dDjuZxM1DrmqSblP2Adf91oyVbF3flYoHTOG1YqX06+7x/AKg+bqSA14YZLBMfQENPYn
x3OL1JMH35HyTV/C4yCnaipot3y1u9cIP/LVofmTvn5Gqjy27Vbg7ll9yACZsmvDH9dfJn28xW5E
qCGV7jD41iLp+F15deefAylB3co6ccZ40gQJ1lkawhhVWxpPmACu48Z7JOPC73aulbLGwOR/wRn+
QcqecrYNf/xirLd9yCrDnvcjXFQV9gKEBUCH4PzunFwhw0j9WEenvmLCA7X+HOO+hd9GYBhKSSt2
L9qt/zQT8Br5Msk0u7x4umXGyyJYWR02sPcGFp2jNEvU3wF035pN+qyi9bm80xEFkam6G7C2zP28
iBaLno2zzLuPxm7FFiVQVcun3yZlyz8QwbIpFH3SDy+Yy3GMX+Ww1RbkMn2186wRR6jVbSNqe9B6
iW5c6AMDcvEbVasYnrKUneKUOThJw1EodvnOwWFAOlpzQ2b7VteaL58S7p2E4SS3RZt8CxMH16ga
ibKNpBpqz9wUCyywJWjIFBgl4XGTaEeLuMRP2McnvaMf1E2joEFYe6iT6ZuTNAKZdp78JwqxeaSu
vSb4FVK0mxVsS6BVfsRcTRrscGy7LqgAR+Z2ttK/iiuolAOuh97gxTCIp7RTJOKzlhncDWMDKg5r
9ax5ukjHpQv0IYPfCquwFoaKQ8Qf/bDYlTlcbeOCkiuOOXpbIzJsRMzgQsVd5KTy3Dwbr+locLcW
YdRB3I/VtpVLluF+nh1LIHrt9gLU2eD7i4qItmJ+BmYiHzr0wGc0Y8oxyhKcLbAzdzxOC0v3gvKY
Ehy0OGKNs43HgeV4xopqjxcFZSSLn8apZAKdwkta06izqvzYPmPkMH15Nlmj62RjPGzl1cBXCxuo
Sx8LFh9NBSYcUr/Enb1j8wgknRsBrwyRmDC+E3LYqCtB1GaVZPhySEjkiCx0EQUA9dn/GV4myQyv
NOyV6q8XkoBskhTOupr6klfjoVPv5dbF/ZT7VLdqwwTQsYssivazphmQxHWbFEFIwMF0f/oD0I/p
ROQWhP9D1Md2edpxZzMPIBOUJ0YGJUTSaWTve1RJGHHJJZN4JHn7DLRPIP1czGbQ60W++w7g6EHR
/FtjDuaK5DPYwtq2bPXmrqNFsw8KiEJwbGEfIZ3odpDq/7FkWT/QPnwZMk8xrPcCtqfKs63OgspJ
cQ7YEHiG0SzIZiLRF0q4mb/w/0DEho4GMN4ALLLKIVXgnsNLeiKLTXpVjiM4YVEcvaodx5DV01C+
trngJbXASozNYnOGJS2GCMut/38nLyrLyHEdtG9D1noyc3wW6Cv0h2Elsnml8byTQhySd9bn7rcS
6Ro9mKN7F7OVnSU/Ho0NSwnntiRmfpDIBk3Qjag78cbwcP9EnC1VKx16/zQAG0atbXd80f5P/8Rc
FNzaleS1XQ82hS00urk/ARZdZn5hwJlob8g7Hvmkn29yCUNfo5ZsC1szT//UoGl7AA/m+oncUgDc
hjHkZLZo/D1yw9DRNwT4Kh00NlyCqEvRc+BTGuxnKsnpvKzoE8/gYa0M+Esf7PgrrrDLRfgwzkz1
tqITQTMXxe1raj0wxwS4Ij/9Cq76/44fyRwYnv4ZRActWMIG72pFE7ell258QIyI3dzvY/4tZj3B
JKMtf5+5oiu6tkGDgY9T7iJ1BxhAfQkVQeEV4GpQilAAHkfEaVBpZ3AoYWKKiWAMRIVJdT/d4drH
lQFR9E6SgB7icXKK6DYLH4mt3jALb0gUQHR3rv1RXn7FCT7yrDx5wAl0Bfg+TalrzCVUAG3Svp3I
L6+PFdwRIT+uAuwDiJgp0QMQjUAyRadKqXdrTB+Wd4mIMKz/zs3svqmaZ0951A7lem3+N6HOUh2Z
1fX0uxox0on8PRVerSsx5D4p2zTkFof+gjLC/puy7lhFYMGe1VQcJu6zvrhE0thmZZyEk+pd9GFe
RxwySVROuKpE7GwA2keumeuJ2GrxwJER+tY1rsti2tVZq29hNwIKMIHl9oOhAmgFxroVJH026UJW
pfPCh8YqJNH+Ah5FYobGNmW/qrMpSGb2KMB1gMToWABybgki64xm5o/at1zY6Te8R6X7EPEmOskK
TQImu4JA0tec1iJmLieSDZugB8ha2G88hgDqnD/zOIWcu9uRbfl06mmMG/2IgCEeeKZl3hs1jgsX
PqO+2510MOQUR9pF3pXXQKo5CohGMhYvF5owrzQ8OdYebwpTZHSKFh+lEBJtiNQw5sYCDGcWC/it
UZoGX1MbSe/aw3P620Vs0kZshAWQqbHZY0SCiEQtdEhe8gESHk86GxM3XVyWI4Rovf8/sjojZqyq
OuLLpJnli7kWXD7tHnrg9VkKr3GmH1vpMO+b8E52Gc3s8D+NUwWOaDWj6wEflAadekOCzr8K1nFr
Gr0B9AiYhCVUXqybzzt/RckYVmUSOY+sAlx7wjjcPnldhJyi3c9CzdLA88jVrdQDlafCzZ51AMoR
tfex/rbJ7ARpNYQ+PEmQqiCldZY9FYCj5asSDLp35sQvv2OBrgBDVxVbvTS8Bg2vyeztZayBFx2C
1dFd+5Hl3qi4285YHEwKrCjDhze2xNuPnuFW8iQj+m8UECYu6R8+XU1llxJCspH5AfsZQutVlyc8
eri5E+Wpf3Hi+flLSxQEsOFsbjj341Y5GAnCpLooqm6+w/dM1USWvPcSNDE4NmYJ60lG12vl/m9x
ybD6Mbgfmuf7O3LUOr+PLF1X0YCB78bLVnv0mAJoLFGrpwPvk41oaYCpDVMIgCKzD+hjNFvBaKs8
TMyBi4CNK/liK5x53rfr6cT7k7Pypux4twjaKEJek6zansBLCKurz9eUnZjglsmE4D/1NRXExAvW
2NPH992HTcZbmGPrDROxVNS37fO2zkfngAo+arn1pcoahcbrVzqHXdRnf4qQ0jL24klbwE6MEmcX
XAOOFbCrOXBd4WCms0SF6buidVjDTtdSKtVjPUM8/9EkVtzsxBcJtnkXI2gZ/8YG7cbiF9W7ngqs
aLFdQMjJLpt9a2azCN6bkp9R8WU0qj3CCdEo74EwsNOknCwUEMCy1Xrnubn6HFBHUQg7O7cJnF04
GxXLMUoqlovSexfntnGO/EtoejRGpyNZdrf0ACZ09ICPKAGVm4oVoSnsP8aEFt111TBVkZE+MF+8
yd+XC3eadGARZje8BViYRe2i890k4S3dQZBzuZqQuXVfu9XTsaw7EinAk5QEg7wXU5eVkjX1ZEOi
knbI9aF63SF6WTfYIPFAqpFN95J90b2tDf2ZF8h1a0t4AVc3rmpxSJ5AerO4lBcfDSCdv2YOw4Lk
/NAcPfvRjBqWlgvQPtovyLCQn3E8OnsyxHfmThVZumedklDbCeehx3Ig6QVM41uAJd3jlL+bXNE2
FjM3B3/TQdSr3uXlwLLunt2szMbwtT4zOvMifoH39QnyUcl4+KN81vxjMGmgpoASDZTlhFyCBXhO
pisO+cJV8NW5EMLbZnMHL/Aop0UmBtgF8sJSYcuEWKGu09CwYqnGSDjQDhucjfhSuV49E9+0Y17P
KfXb8qs3NTnzqUGNXHqT6jn6oxhcWPBH+5rYWWai6pB4P9JTqDJNmM4ajf7x2MC+7zCdiv11xqdg
7PVAMAFsS0NXYIe5EF+Xtd+8AXgnepsrSpoeOmDjNjwhlfFnsfHw9W2WLAuTrIWlzGwB7v/mPdT0
zK89b3lYhwllaft/Lw0kkl58d9s4vYiI88WZYJ8xV/EXVtBqn0OXiWwP9H11IzaH9D7cskOBOIZv
RUNYck1khESSKCjaxU5Z7OlWbBfowkF1J1hawPRMtcIPx+2sbvUNW/TKbj8o4vnjN84cfmIXgnqH
81wvbCsHbGcpMh91+B6jGpMTVao1L60kRujzJcYCnIPLALZ61ObNTCyFf6l1iHD6PxglQ2iPXD6V
1H596rfYogB+gcPn4h5PTkjyGjdWMcq2DIuKwile7wsmbrO9TXsEJVE0eg72ZjwoVXD2Gil4mmzk
E2b4rHrkXUb2oGPrfHEji/zRuIbmXN3PCDGmNLBoPiU1Qv2SBFGK6OfJJqKusZUu5N3RbKKROZcM
vsJ4GV2Fen5RyoTj+n9981AklpQusXmQfErGaPaWLjZw3EmQ2JkQnqSLB/9bqqEhleWzCppbbltv
jr17XnMfobgx1iQWAogvO4uwmIfyVLuKFPXu99kdnzqMJXN7PB1J0XRjxV9WMHKh5Yka3sL12TCB
mdRRsNwBDgrS8mHuzGYHUaTclsnk9+L3uNUwaPyXxs73K2Pdozi/PrJQf1zUZPgQjESzbxKnlJRy
SBVmCIhsA6LIVtBug2tE96TLivtICnUcpAylovn8YwvY0084l8803kTHWNxvQsH+00+0ejR9j6h5
kgEdVHgwmpG1PvwCxZg7NPCZUw1UpiwnGvgkZ0tpbxNbYF9NH7x3Bu1B64vimsv4+6qDkFot9ypq
Ntl1xqm9lw99KKcqI8e4EjaAIpGLPEaz6iRbOruFq+auZuNHl/BviyZa
`protect end_protected
