`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nxg4I/GiciNsFTX+s2NXWH8uhH+SxHYkrfgaUDVgwOkAdgixTuWeIwrIJ8nb6IZyVDCJTJz1GOnu
KVT6g090Qw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dtu2xDN4251ZI15yhvQNFpogdlJrqrJb3b7Zh4jryzhQEmZ7PWDTWvxYzP+adlS4Djpm1Hhh2QN0
5ImkDqzKGV9e9toYvogqk2JYKheD3d4fSb8Lwswnhh1qoGDYvYTMAm+ZokNn9gpEnbqixYmMrfKo
xMj5Yq2I8FmYEoP3lJk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iGRrx4eYWh0u0meFsC6T9928o9OKqE4shhYxaPjRXZFuSxj8J9GTuOWOndzAWHmUI0IOfVykNH+j
dHmz/+npD04tKjRvbj+1sEgngcQg451W0kRWVcG5YoubaqGM2wKgVJ8fshcKwS67LYOtch8nVNBC
o7bT/+Bj5I/ssYWDoKuI+gOqQ5rPnkPPk5NcMHDTFNUE/NqTYQ3+x9h/WCLZe31k6ITFp1bX6jYn
C/xnvCXs71lHo/RbghHI+t+iUCC3RqvDB5agJfrQOPVmMRSSWkNBJJXrQ7R0LDti2WacwXS0cWDo
XGt7AMkN2VyQ5m6Yrr8yiEMdBC2lf/KhidR1/A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zktREDzfH2/9y5/1C0iceh02VBBzhG0sy9mXKKJllrATqsxuY6P0/MQL4OXVLODfqmVtQK1vfpuR
r2BalOcvNSXGNJSMaC7yf0xodFkiNhsUG0DN/Tub/N7xl2gYYzZP4gnVpIzhZwtdhqPLLmA50h34
qSNZTkINLYCR7B1utwM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oyXwtsFZPQK7VNM9XAoaSGfUOt4TTHVcE6WcSAjq278Zxq6H+Lq8s1j5E+JFCP9HrMy9hnBrzvtl
+LGQd57r2iEkNvGN+ua649Bjd2AXjYxI7uiAE6eGQp6GelIb6ElZMMfFrBLM4eUbSACWdzColWOR
xCypk+m+UxlJX+G4LScGrn2Nbpllxf8poFz8nwbYNY3oX+5dJuRR1minN1O1U9GCP7fR6cqFVCaj
L6xeyN0bK4MmRLqsCybq5QWNKD0p7RivZPi1wvMTmCGe+RCd7ieX0b/zFX8VQ1QkEqyQqnh0BX7G
sVbhtZJkHBWk3I2wpOlryGLZdr0kOcGPZ8qDXw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3280)
`protect data_block
zpXzm2za1ZRtAcd2O4XX0n5V3P6PSR5glSylPkE2oswdfooyMtH3q5P78+6FyWhUkrF4sklrZGmq
wmmvXkwCxOGSpRkYkCXdy8WJ4fzIgHhWxy0oUMA0J2Hnr5yKZEiMN+PQsQLuuEPn7PRT4+gSBvye
IIvFOf0DaRxbMzLhxZwLO/6Io8mR96RtmMlqb7chtO5g6+K76UjzAU7glXfqOUsAHHwC4YQk9tcH
W726wJjaboT/An74Mgj2jgQp8xsXIuEn1XikV3iPXe2Z4ocWyxExCs0OSykibQY3fr3Or3KncCXU
xsyCM1Ap9rUgk3u/RCoFsaLGRiy/dSXkPyLgGQRoZZxOHU8l19/o493xaknLKtdEkuSDCMHQOPsc
zyeowhp1AgUQ4ZXDQlVvFyHn258B3mBc4bNZOQUk0qf/8NaAm3tXEjMD/vUMGEFHQpsWBhZ4MeuV
9TqwWnv5WXFd2ON8KQ3bZjw0Sg0qsakJFob9YGuHlvTfVJMYheeEjhHrDrKCc7Mgz55mJK6anLd4
xAH+QJ8z579hmmR1Rh083HhPl1tOht2+2gscK2J4FeS0t2NVWlxbGee7WEz2j7S0zHBy0H11hd31
G39IGVfjuw6Cf/gUQQ4fmLCeTj+YgvqcMYSBnN+PZO9/4WYidwmEGJdSkWGWqs/VqxJ3YmVUVx5l
Oss4V+G2i+2zDtbPfpGQF8uqA+r8byaeyN5WP4RL/rZ9HZiW8KoVwTYNhHU7gWaefgLbEMH6VMJo
luJpH4L0/m/6Dh2Cph7DDgKAOZKjYWdL50laYmZyUETvNf/nS1W/IPpFZPUH3ZCrbrjoS+zLI4ap
TWWw28aLZEbhdtAte2v0+3E1GwcW3fsvqb4hDnhDSjm/vBQnIdHtNaTZ7FnHwH9hCDDXCs/aggMz
uGf6pBz+qfus7Q5Eu7QGWc3nESO8Wl74FjwqHiwSNa+GqxyedN4BgrG6cb61YJvGyKjhNi5ONolg
5iXh9tt/Hcu9lpDnYWEpUCpdibm0iW79vyd3xl4JYcbi0tVA0OnIAPIKvWsX0kyt81zXi8A4Ftyz
jM/5/EEndFTR0j6Mh+DUhLrxZpLRtL8kTTbqhipGKPjOhlB8l7tw0Xc2nRbcRGwSp8Te90yNBSJy
3TqbGfm+lc37g4MpE78vi07/W7gNtJsIY4wq9WXFWxogKkLx2aaaAjN5hIaaG2B++Hvs93D/lcYr
9l/INncl2j7FRt5n5WIQrNPnFVwE93Ed9U2SYhu0Btxvkfw1kyou7tODzzYdnhVzN+KZe11LYp7J
LGsnQDD9tqXzVMu/jNrwGvFhSRaouh/gkE4EWuO4C8hTAzK0FurXuPFgvK9Di8PyAAgkD7HF7EWB
BDSl9mvmkaMyUt2V1sH1W56cwQ6LWsgIVuBWL/jx9X8cC2hARIiq1lOtCPNWUd2K6jKl+xvd8ccs
EIzWjcsHd6hunu2laaoNeLG5FGwvW1HxbJRIOZ89EEht+BSnxTt4fP/J8+TYBs2//9OkZRIAsHxC
HxON0rymhKrplACVZMnoz36OJ0qY6YbHwxI1/CEQFx6n96mzP6e1Q8SDsaCAxvn55Otj3aAzq0I2
wOZ/Wl3CBgXC9HC2jezLjTsb/TGoV8qU+jxAqfySs+TqzLVqhyS+Px3Bv/2cbaHlrqSi06z5PsHD
ktkEizlxkX19q3YtwdJXIoEEZVOJzVurRbvrEGB7H61XqwvrvZ8N6towv0AM7lR+ZkVtnGXYkoSU
DO/Y0C779HT9f7tUfLmEbDfJDgJtj45CfX7qJJg+jZHOmng8uwCoZ0S1c6NWHPsQEs9Z7aQbCqc1
Yk1ZMO5BdquuSvCJ9xMFhbktFHlQd5Qg/jVcuxxG+Oi51ImUgXEqlju95RVnoGLjc5hhCNxpPsU4
Y/uDE5uhiwAIlNUeweqtPvACaR8RfOg5D+gOuVOavi96D2cOKFsarjSMqSEdJmeQKcK1y1RF1GBL
QTmRDvjWKnRD4QeA14/5dkFGoW4PFmUMruSmrlVZSRZEFyWRp1qhzips9zXvyIK1Z5PiGWD5bMg+
qA88OhU9rJkMZAKYMg0Czew2uCISxZHzVx9HncRbNURIfsb/zBM2yJFVIvYBqxal0EdMFE9gA3y/
P4Cy+iI9qu1lZqlq75Z8Xjm/e1HWG1M0T5e8bLLxc2mFUtIvXrby7USMshH4u6WjOhW6hQDBZnK2
qzB5rB+n8MysqN7lFAES0+b4pNpeP4xy162V6rENAMPW7rkWhWsYv+X8lIa4AcbIJQ5ntK9t6USI
6JdzlUb78KdntmhD/lE5QYOA6vV9W0AhwxK4bZif1Zh6iieJnin4KyJLP0RrgeRwzy9CQMaQ6zbY
ddZ68nII0BDnnyvangAftCM7l96jkQM8zAF990t/7YgLvoDnUs87Pk2pnqDMdTFy5zb5anJWtqFo
IsJ+VfEHje37LV2uNgJ4bI8LuWHH03ia9Ne9Gqu2mmw16gm7+7AMqOiTyU0xXWeY6wAwpwvKAK1g
eA88md7SjXvMWHlfebcjRq+twU0V7r3oztzwcclTpwEm8WPecXt6wgffkYTcMLBmjbK6UoBfE/Oa
uPUnBm8t2GtacgZx2o1LkrQP8Ey6VRP9uQqDq9Q7JcKKh776eWoTuR5jclwkD8p+wMyequ/JfyC9
8aY5MWkzC31iafOfkRUfkkPYYzMPmXotDGFwNOYv2EjKAMbhr4nV7cbqc+Y4Ccc8tRfcBzlwoQ/h
Gk5t6roNaktrcB/sFcb42S/8OF7pMKkPt6mp/9rIGC6P669vbH5U7cJtWsuONkitn5ptxVAq1kjg
Ux80i4vsOZFJhRrpn5SkRzjFM+wQqRrhqPTwTujMq5f75Vm/GeB60P4gF82ytVel1vjG265Ykx88
fgsUbt+muAkh2n5g3gQ7bH49VQrfz3nDeS4V5t+/u+VsDeNSGxlZvpGTPSREU4CPM7s59+pYur6f
jbLpPLfOnCnsTpirZm5Bf7zfEjBYVi6l79WEzJXxxAvyLiykqYoSqZgR6c8bKl0Ic4UrIRxBpVx2
DX3SDmoGCBHWF56BtsAf+t/EZijiyPbAPWtY8uR6b7RIFq4pOs0Wfnwsnnu0dM+dQh4fIMKupHyb
jwDtCyzbGrJa70Z8oLzLzsNoLk6fRz5GNy8cUzgzHe/0HHUFpLTNRsHw9sAbArvT4CZGHSj3/H9R
1smmD9KBZloLpgagmH1du4daZKBRDTbTozTo70DdvJljC+mH9kpqpX3+68jEnlm8ryBJd+Totg8u
nfuBgg/lEbwCkK8EnxidkYGpETRu4IbIYsDNMzleyiEls6AtGHCN6Z7AN6mEuBOAFs3lOyQxNtA9
yFKjGR6le21WiPMeuh4Dg9z6G2El9rEPaI/t+J1e51DlCO4pD8WdgQvPRBoBR5DBENwxYgWvfrFw
bidixca7zjFBO/0apFVSLlgaLLO0N7DcbXOFUlJlx7j+ZnNzvKlSjbKazCe7R7QU14uaQVYT3sGL
/DJAwRCeY17mubJcHqlssWGscH+9mpzGqdSrZAzb3KJ3EHXry1IgzkZYNgvVfywC79LyH40TMj0z
++Hox5DOMCY54D9P+Zh7EDHx87TdHn4yd8KkqqmbigISsAtQj4hQ5N8MH/sEisqtma4vwSevOg1O
DyQK1FszVtcBaZsKFRxWdbv1ZHZVsvh8gebbyCFJTCnPAhPYigvFrxwGRqC46teaLLPq2pB8aguN
A+qmfnhyNQ62pVKGwJ82XE4c8nHbGCrdlB4uKi3HbbGRnLFDN/tz0T4iNpJCyYNi0tCqm6utQ8vI
674ZIPJ4fp39Sbrvd39VvyiEdavytg95foqhwoyUIN1IWJXRsm267HATzeeDM64eEmvgpCTwRpnv
X7LW5YE4whYPtA83YQhrhh29+VCAHHW15ECUn3wJYQ5/V6qd+eEE7R/v7wbzjPBMoG37nRNk+A1s
xDuybfKg6vrQTdsbu0QoHdbL31qR0cnZg2q0OTGulKlpNf7Y75kHFFOZGxyhJTvojE2z/YXzJnAL
MKaSYHjAWJSxBycaWgPKy4DcwD8gDPSZi/cZ3OM9165wvw/toAeEuaNygpPY9vP5809qtBnCVJKE
Gqb64v6Q95fDPh4pFuSi3vGSNKc2O7jPIjptbRgN+X5LdObZxYrutX3x2ry8nbUBeFRK8teRhqgH
SaAO/XHzZ3niwYeL9DHLvR3a9TO9wDXf4KQbONTmX3gq7pIdiAUpbqkqjEf9a1wdyR46sd/iX9hh
J+0C6lIjBsB/mEXcexxwqrzGZAKycUJG5L5gB4c/TG7dLAajrgTsZnhPFeEnpcx+MLlBlXemueZs
Up7nF1My+pWNob+EKIUMdtKmm6fHg8MLRAV+9LVMMg==
`protect end_protected
