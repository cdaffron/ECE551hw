`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
egyvtHl2SqiIWuxYRtM/Gf1OxulJTylmJWSdxw6I5J+YJrFwSPwBqWKNZQiNipAj9STMHt33rdGT
viZEOrKlRg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m6XnLZ2VlyEB3m09l1entatKXbnODi/jkkJtmibwwsB/dYhno8zilP5FxIwBh/7nIsfGdCRzSZIk
y+sHlzpJTE4FgSvf9CHgiHl543w8fw71BlWzZW6dmrZGCAy6JOlYaOmr+B9wYhO25gNt7myui9i4
LAURT8TQSFk7nWsKDv4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KtnNab/js7Q/j9k+oUY9x9R763dGpU6xKQj5fDSXi5pLxbQN4wnNUNbIe5JwbMhncI2FRBhyQCTX
gKAvMmLOilRia2ps7j5auCRGE5y3N546QfrxNPhPwWjF05kRSkH5HFfQ7PsiC6mAFqDevCfcg9Fh
fQ8NI4ZfxnSYDOS6/kNZFSStfLeO3IAy7zOTyV+iV6cT67hXxSjsmVL2KlPF+K/XHBQBBgUofFAi
N7yoHotOeUG631i0i/Rn2bej/eB3eiQTCeeEN6OT4pVABO6t9C1q9IIR3bXapYlyp55yFV1hz5yu
xF73S42aQTaCXolafQ7KrzbNIc3m5VWrefFBsg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tenuQ4VBb5Ey55hWgdiBhVbWwGDdd03QKQPXkJjcGxQiag90ECKQ5ySzzjNGGK3lZQQH9AmtByQN
7K6JB7Gf5Jr3Pr6uFuSjvORpVFi27TialCaOinGJAbcrzyzsB1E1rPOKHt4Jj/eFX3AiMle2XxPh
TbFBIT/1boy+JgAR0Uw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pgu6E1ZK3SP0aZk0yKu8wW4HqYUySdFkNak/SD4wI6P+6bSpP0N8qAqhnObwKJCFHVusB8I+kKz/
JmURjLknpLA9mQg+S3o/LLoZfUUod3+9YF8+grk1jrGJQnpRCK8E6ZcHiU6E3eXx0miGDl7Oz/JN
PJaCAe1yof7XnpzawQ4IiPeKQLRlV3/I74bFSx6OuKQIUi6m9DHqI+rM/HGaMx/6Bgrodv2DDlMk
Rxuo0OhLBPlGveCFahobEX9cwPZ4aJrTdRNE8EFvRPVS9xxvkwvE5eJBcOVGtGYFqg0GEGq3iWHV
58Hh2ezW6wucaGnIi2UNnlDUGjWfka9Fx3bsIg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5856)
`protect data_block
EMfZp4+Tcz7yBYvLS4kYGcuvhOkoh1bicpBUds01nJvzYZIH/wZeyVE2HXl9gomrZbWtLHt8Y0mA
ER6WJXmgbSFtZ+wGRxKrduHOHHlZW4BNOayM8UiWeYCXJC0CWdJL8/mehN+uzY658jAhOotxWabF
auRbzvT+fVVfc1J1YLpqUnWK6gSqy6J69wH2WX5fvRC0JkufBejjR217IzHv9459OQEgOMRPdv3y
KkubM0JnB9PYAORXI9Nlwdyw4zLcCEo6DKmx28/5+fAb7d73FIO9RjHzgeTztdyn80GYh9fmUY8S
QHQJqKrCHXgpR5RYnfo/i54NWhOD7SzPgNNg0mfLMk4acHP04ppsnwZGxQlGZLE9IZL6LdtflBYX
NrsWVkGcZYFVKuB4t+g7zO3ktK33qEEzd2jQB9DAhy/DvB/oIcSNYLGuiskOCv+QozdorncjpsP5
9uxDZMIPVoV6cutfv75ET6RGAbImExQxycw0mbV1RQd56O9CwADKs2SDyoTMMqvRz3KBgn0LnrNZ
RQANzI/6RoKxHFem9shUrnlCESPBqib4/EXKadpu1qzzS2znDIUs5TV3LyYpBfa6vZWcqseSMlbX
IySOwasOL/ZcVaVBAzO/yOLDElpknRirxP2AVRdpo7Opkx4emnNweAmYzz8WhfoQkwdyEvIsxJkL
s77yhieP6Fj7l9aoi+I4VqKTb8g8I07wxWktkPjPcndnmXmQnG6kCMYcEe0aa6jzIpB/qHbpALFd
6Q0sC1jbagP8nwO7QzDExQQLwfbwUMYJIgc34oaOKJoajF7EtDFZgRQIC8PN0NgbMMMPA5wIQdXP
b5Ak2zVZQqA+h3qzwZ+AAjsdh4yYCUGH6hgzsfzhwSKBodSwK+jIBTlW0O/i/1ozBEr9HNSPC2CG
YAEMZcs2JymDsLcFhtWxKWMjQM9oa8yk0GrCjrjejIK4doyhcBdb9NeXvBkRFhXtJV2K2Ock8nv7
keZxTffMGTT+OZv1TJYDYK/bgkwbOlMWekBTShtJWGSTi2EWGWvHrQDvu3GvbvfS6ZxzxkzlboFQ
8S7ui5MyTylTCtsNhFG/ABR2nU7MRdjU9FwCL8uNPkgpFZLcRBYGW1/Rr1Y1OAAKQkYd2QKjrxD4
Z9b9DKPOW6u3DPM73J9W4eXG/dcluyvWtCTkdhNGcXYHQjWa3WbQxUfPJRjVjWl1yKnbnyQ2GpNL
01gFTzGkzSJ2NLN1T9feRzsCahWhsvP29302+NhS9tRQAUgeNYEDBlOBgz762xWhDYqPI8yzz66J
F3ZXPr5AjXwlev3Lx+es9XujxzyY36j37hTHVyymniJZ0QKM9+Uxaf2S3trJhqS0c45m+6hvxSF+
eW22YlA6+lAynH0JDRzeg3C/PxVY7UqLHkyLeZ8g77xaMa+CjDF8Vhbpr7MwY9q3MxV0LSRVT0A6
gtwPm4aurRpUz+YeMiAPQa+CIB1RrPqXA+SxioKm4ykIDjNlESqd5O7nEu2DrNrXHuLtYdGS/BaS
pW3k8k3h7w4fyYodmelAR8BjBx7E4rfXDDqzHAAfT8SMhJaTz9yFAqGOSUVwqVh99aUQU3PQgIG7
Ji3szaYC5GHg5lUzCt2vTwFfPNX0jGmN0f4l0UwXbJOLskydu6r201JCGvi5xrJYiSbCD54qeWnH
EQkoa1TNGlRpDtr5RcQ6RYbi8kQy+q+pSsvWTKwS8fJSqTRkeAfUNBoSI/6SSSuTjhLxc/puWCh6
L4soGGXzaniMH+fJtESuseMjb4Hj6VqSDRcAx6Kck8KsXXGrWMp6XcL7a5gnkysFpQ0wUCQKznLj
6moKTwtf7F/B8tP8DPX3AA5iqvXgjAJy9GRjzHqPFSID976WBnytf+NK5zohde+ugR1x0+6t9lJN
KW49KPx4RETz7Q4I2fmnO4Gr/sCYEImSScefeevE0BexNAiAp+vrJGG1pyk76GC1a4LPrFAg16HJ
IFoHTboZGoTjrUFXDrd3e2xtGDnhBYFiwFwiy2b1RsEdZA7L6bk+zgJuvdY1Y1LmwEcxLjhgD76M
SW/KH8a4jA1egNYWH9Q46f6DOUznSJJ58ltGUYymrJ70+DLVbvn+ys+xGC4CdTTN8kh9+YN2+35l
XmbLyYejrrOxjZJHw+/DER/aznhYQV10GZ1pWwzf2Do48Bct3yUDRrFjOa07w/E4Pkp0tbM1886D
3HFPOhlbHJ1MzEG4CZpweaEWRqFjT/AO2TXOhwhvzT8opUEa2vrPjaQjC6m9UJDmbVBiIXZ3G1UC
ld3qS5acIZ0kvXPC99XS5SabI2e+0J1rbwStvutSQ0c4Hcsqdb9OQXqrDZtPLDpFWnGxbYHGl7nb
IW1lF8x0baZYWKCFUT93gVMJ79Ya4f7LFvt50/sMp0z5iY15sTpvoEbc4Nh5egMscHRzJd3HGFBn
DFBaymF8gUGN5BRpcNkCk2iGw0aFeCZLV/4hTuVzLvZlqcRNdFybkMQED4O+Nq25q+rV0mOTLUCc
3/KKwkngjSOG0EsuV9yppXomBAj34H4SViWtrpeZDBWIIATNRjpMJgDZiCTS/dCSyOsatEBYaGeP
Ech8F8i02a0vKABIYuLo6p5jnSXDhnCCuDP2IRTUCDxtR4KXMUcwFuzRuanD0Yjk30blpFxF9fP+
eJGAFDwckp0vEY3iknrqeX4ZJghDHbGJbGpTs8hQBZMIWUZhHxdQuWUYO5JfsxbyqrYB4XmdZAvL
MY3pL4ujmySqkd8d+3WoUt5d9ti37X4awvRIge+s+rIYiDTaydrVPvx1Tqho9Q96CRY8YISucrNm
F/Iqgn3AlWfPID0sEJe74dXpw7iSSdMwAoX6r6ykDXcTw/58BZD2CA5BtMmc9i6gsM4dwgjI/2/R
lPSq7Cr0m+FSsPmDPyULnEJRqu4QJA5bcDIfO0IHt5r7UPE8uLtd4O3yvEWBqMU0b6Lnbn9kOWrX
HCyG/mC1n72CkoEZZeuv0ak1TxL+N9PByqbztaF8RRk7Va32HjdktZgmY89Z0uwziCZF3Z0TkyIW
rddk50b2dhSlSxgaC78dWF2wbdhNLp6a9KDhMbV7JqiCnaI+7vwwrzFHodu/D+h2g1D2kXqIfb0K
7XeBCBpsI94wZ8aaZTW4S3OIbpOUMqnAT6nM76yE4TwROa0DNszBsgND8KdDs/lbXb7Sr8Qc1NQU
+B0xxK5iYJVWx3orQQXGLSzhjf4Z4JCYo3JxmaD+jF25Q7ewBVZQK0STDkbuIUXSNsr85hUYXhG/
j3L5xor4gEnabKyix91E+ArrulQIUyIQvLE5YZS+uHWj+EVyW8B01rkVTGwJz4rCCoaUH4Sm8yYb
39vS7XYTasrviB4MtqsqeMyK673S2z3fsMxLuLRBMkagUQF1smKOwHiFCbgYzVTRhqQObOC4INuk
WSoQHdYONR9BMJU46Oe2CQoeHvpaAtxmvyfxAdYJP9mh0eq3QCait//Ff5dF2HrqHl4rEebgUZDv
/cVQDQZIiBdZiffHEO0d5VmfOAfa335fD5/lTHj6U1xqaOmu+ZFqAR15SBv0mW0LsHxPwjCzEnFf
WI1YCD2ctuvtlb8/EPwlIVv+x2Ey4O1ZyBgRrot5vvGlaydojBmKcp84DOCQo7RIswLAhWxK3pdH
T92kv5mZZu5xJh+BowmHcsLGzTuwVfa6Ur4p0JRYNoVBrjNUrxPCbB3wt/dz0RY38tDGpIUevJHg
K6ePXT6W8tPpy8tugA444PjMOf3I779dzyUlK77ghP8ECS31XKz2TiW4odJI25lBKjqi4n5ErxKY
CqLt6/dVCuUaFUZU/uRC5E21QdALmBzRho022WVqpF1LU+ZArQlvZt0ZGrG0YJ0so6gKrCv5aDya
4Vb7FHvTBTv0rTaHHvHzGvWkPWHmaYJWC5fx4eVFw0f0I53nKcY7K4ODvhfJ9pBha5XQrETkUlkU
SoIZweDrKP0vM7WcBzudKhYfe/IhcyHMT6sKUWWJPzLfaZNiVCnN1OkKaaTHUXLR6rSUcwgSmO2o
JQKnLDYhI6hHmcU49KI+htt5i2qZw4AwOdz7Dg0pG6Ob0EQYRILdLbLHffEVvaGWsKufW9YWp0Cy
ZO9HusPHTxaiFWpH5inGLRyefpzS+2xZUVl3KlSet+lGRH97OjPkXzomW2uW1x0Zsbk7/VJbor4r
Gz6fA1IJEW+CByLa+0jmPqrfedGyI+NS2zCwCmArHefVmUiXl/sZpkWOBRsla5MpJCwK0MFsMIKn
O2nD7tUFRdUVCyYckVaPi+zk7Xb3hva8UKAKLIZUWxnl5qaieXCv0fiHtmOLUV1eEoIyC3E93HMU
qJN6u4/0B/X1MnhLHmuy3JGiZzCihETTa8HzsPxJWIyaOJOTZs9VA6KsrMtvZK3xv2oY+Pjvod3M
49+cZiZ6sR8AXShGIdQxk7/i5bRbOO4EwXmQy72SwsLrPBmm7cBHPqn20P2oadRw6TyVrvphocdV
B4WSjjgRErH5tMYILEaSXGYfBDcxggldKhR+1BTr8HMerwQZ1ZecoCiW5Fo4zDTawfBO6E8T6a/Y
v9/MDEu3MhzMiV+p/u8mW4759DARdhX9ZBnuP1WhtfF+Cg6Lw2iuHOpAS44u0nEPgXgkR3ojIXXy
CW8m91x6US7E39lRDtCr95f9n6/AE0ZsN4W1CVwsx3xBMRsiTk1Fl0K3rpOSFkkuFOOSfF1BQ52N
HgGtuxS6qUnWHnUt0c+xCB+R+MsCFSKfHI5yfWAltfq2NEbwQcU4qUpRIzvwB3CtpX5+qmvn3wGB
vSwp/DRUGrzGFeq36/pvOvJdyKsxVmM4tTTOHP8L6dgC+HD2PvunZsb9Wvz1FQFEwlem/nMNUkbD
XiyuutbUcq3+YKP6aeHgiYnVLL9ng5I0eP3+xC06/ks9V+H5JerUAeVXhpk673+Zl8k1WwXAdRuk
KpX2bDZNKTlJbuG9Sz6ELp09YbWS9pmrPWy4C0EmCbIhSEVO4l5ia3BPnS3ox1eXVsH+gy08lNzH
QqEEUUFvNedWK7vENdsMW4osq2GpGCRIn4IdH216mslfKhsLBmjI/BN1m+UQ3Qx6G1e3LkaA25VA
afa+H39MprcQAPo6p1AbiU2gsHZHiRS6QTvrYLL8Bze5xYqfSUU1W8Wa5i+pX+VeNEqOC3wH8gJY
AYpgfgQ3u9Zkoi2veQHd6ReF1xJBRRnBPiWK1l7/+LC3eVG5MxnTvm3u7d3xYT+Ioa/TIf/AUhve
7phQay+Fwc8kdpzGwQ4CDm8zYBDwH6xbCqmxXMEn9E4YxjkZ6x37ywh6vcKK7QFSWxRY4atWWI+Y
RwAQiKBmwjziGAjVo+M117F2JyfNa0WN0Ow+qalg0wuSdOwbyGKr20IkDP2BaLtWsCc/VkJwZE0w
WsiKcMmK6wkqEllj47tVnBSIjsZ7Wy714W6PjqmM7mkQL4HILEA9vqU91fLowaMyXI8OdqZ7fP1/
Uv2VEIO0V1ZeVluHSf9h24iF3oyQRQD6yQ4VB51RGyrIFi28wUiZZGEvz1QscaydX0LA0ddI/cK/
kaGOzccs5+V763rIy6kQiF7+OWKvzqrQ9B1Jgzn1/3ClxInnRVHEKmzZ5Er3TxnCRG7j87IC//Q6
hXS/RDjshmAi6U0Mmp8BC7ZznXA/WvxCXfEgLnQ2aXVCYJnG8wVN9lvduJCTV2v/fUTt2wviJjH+
OlRj1wzFosSy3RWAtOILc4QYK+3utCUsfeqqKbIxbF/3v2OZj/lq5IuLzxjdGLRO0NyYNEpy2NUL
oLIQoOU4KxY72u1RyWjkCqYDGpVDlSqMx+K/e+wgAuQwmQo2h2n446NQzZD3F54cwMhKxN6VJfvz
f0L8Dx2ylIQxllEVAXaIR25BNjy6XUO9EdnBmiiRVLLZmT7f+cHDzc2RdAAqOPJXCGu0P1nIlWVi
OehHT5qAEp0Fdq2GVBpOL+CEhKDMWOdYvMkRYaTQucxP0rrKDpN7jNFLyGkSbMKT2/ixxoSh/sc7
X0btVsE7n0sMfIpdTjSmr7Ee593mfRnVoE13yrsauTAV2nxXxYb/Mv5q81Mjcg9Cszg/osmv0l71
DzHYb0BoMeAOQLllkqItxSnygmTiBMRNm3tvNwUSVoz9xUk/qOiQTBAxtbicHRJji0mHayoKp2cr
/A/rk39ty0TUFaTkKEkWqmhHZhrqSOHNdkSt4JTpr4Tl5icRnK3cpw78UreznCxBqCLlKffgCw2X
ckD2PzA/4u4rAPIxTCXNcBt0IgrTLX8+dMXbqxs2DqJNeoYV8Hr03m+EX/sj+Afz9DipC0Uf2N0u
KqPV1iPBho8eT3LWoJ+hngohJMyL1VtupnlOFCBK2YsgyZxnqzy8apEc/4e1m31AQybso8HZB4+u
6QQ+7Dw/MZNdbGPo/YWKifhqedm+7eFT/YmOZ2ScoWCv8RafVNudXw+eVsvdcYRrr20QC/lAE7Oh
yrQqYAgLwxq77D944r8XDCnRkZhKQ6mx3XteO1cQgEcXntFkN6ME2+cZ3ENiOSuj3roC1BnB9X/W
VoEy1Ob46XRrjHCzT0mGLDSl+NrBT2M4ovchtOjkRNSQ9aGS4P48M/hdGuFsTK9LElaHj4v/izOp
vykYthfSWOQyrlIx6j6hbG1pfbmWLRWkb1chRZv4Gy3ngviRHaLd6re9QTefqcmuMTP+aqSsaFxt
XgIjO7831fYsbxI3Heba8qw4hM4UU8zcKTSAefJH7DPMK58fN/zJ/5VNb2IOOW0RfqDaENMuAoFV
rboOwH3E/vTwlv4UjiAAHlwEmCmifhwRspTr7walAfoCU1AjmVqnn25eZF/DTpnNuLJqKWyJu03B
QjRbkSl463Wu1Cw7tNU6ISnuocRAmSNl4kGPk9CwQZ1WXYUE7UFxmtt+iNLXhuzgibKGvgP+JDc3
yUH6BEZcASExnk3ZFuBgo2i4Bkwdr6jrUksSkE/1Buk2LfSxsnVhqjgTZ2yDUXnh57RclldLbd8Y
c929HvSfqleLL5/KEEgt9Qsg3Zvw6cMirsNhn+b+l5rok9mon92niviSCuG3T50WDDL4SKlwz3wh
XU6Gmk0DDxz37CCO9vlHY+qVeL1KsiXgpJtmQM8vA13m0i8NlEV9dShQi47p4lrGaL9yFXEFeRQF
gD56e9ik2jSCM7a8bViTTuCRUZj472it4ADikhdhKWo4p6C0iJ5eDBolIkvRHBTHM4nJC80Jcr0e
5v7OWbuyAfbgv39jnsyUH1cUm0Af6kti/dh4afnn4Hv2VuHwe0lusbMFrcPfZQVcO98nmTMJn4Ss
dArbUMDVrgQ+e3wthduviU7KVddeGk3+0PzNuqEUlTI3UO3i1O2e4tL23O5jLKqzEtdeWsffzb+A
RX13XbOjUZ4jIv2MPXu7tjNVp4gmsSXhGVg/GPGlgxREo62TUsPql6j6MlRoTnKUy8GVxMFC4M7p
/09TaUS3id/iSkq0cZ70XWzwW1dct9pe2dgHcuHf6r+iXCB3BhI4luv/R3STsfSR+TRUT9qoAcFE
TZ/nXZtn1M7llMxc8L8kYHBDIhYCgIWBFaoyWqV96RNh5CwfrMVl6Bwnqyu0ETelk9T/6nZs24mW
PH5acVDUIV6TVbp5NGocZQBpd4IHgm/ckexjeojkQUX9xZQvm+Nbo9BkRJOvZd6AVQVcD5OD56Up
LATXDGxI5IEJl+eW5t03QHTrKIDvrEW25urN9GStFcYFKLWxyfjIZMWeol+hPv+nqnXdkv+kkrZA
eiGPbHIHfQ1uunPotLooXexggBWd7TYr/MKMdmyLopf4wYwQU04/o4Eb
`protect end_protected
