`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HDXikpAbEHY3l/y0jXSmh642iwf+6b6cQ/yiuUF7vmPRD90ZwWnt5d9qELk7lFq8k4BpYpJqwQwE
nlqMrDd/Yw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GfKMJiNAYc6aRTFthrb2wKNRxXHTtvEbOCg5qVZrAVxr4a5BZSibT87upq8wszE+BYcCNq0IWiAG
o6x3h/NAYXtYAWIsiU36zP6SNjUInkPqBkS+mEj0lxZiUzcduZPTnLcAmituJRod+tYVfZgsV7W8
2yLpvTomn5Oo47DXz00=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q/OFKwc/06BqfQUaC4cNiF0WA/ms7+RN3L2WIswIciVseFgOKk1bIU8icc8Xl9ouMqAx5ihpaSiX
Z2ai2idOMfgthaFbS1MYPEo/yhJUErDu8tLONreBCl6m6Rks5u46nlzCnnjEWtdPxk7JUtjupIWb
m0KVGKvttJgzE/ieDMz6x3mXQQ7TWagtOaoyGcs+LCOXghcFDQdjxr7Xq9jCKadmArkQAh+uqLOv
eIgFPqJJrv6M183pKza9qIg6hs6NREsh7uzrh79Ctizx6dGLdRK6oh41dmbfCA22R4Joq/8YydCG
7ImT5uf1GNweqlkTSUv0p00w73x/D7JS3pzt6Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ENOA+EZnHLmlJOAc5Xa4o3rWp8AS/mf/PL7gS3zCZYaO/rZXsrOSvJ3DunyCnyim2Hv2jCAoTSYc
wV22JDvYFIsB6YjpaLUUB0Hnu/z23dS6+Vz7URnDius4LRJPBsMkRrhtCiAzIQKbkr1iVfXq+I8O
AytUEdumqhTvZKPECYo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q8ahOfZhRKY3Fc/JT2lfPQD4bMKBANeReJHlWhaxAyPJQISkOJzWLffTQxoGYhuYszF24pW91Esl
O+09cMfZRDBXOaThaW2X0CVcsjEpXpSvocoVl8h7dhkZjf3YMPjSd2eFJ9O1UIuVStYubQX6szRU
hZs7Xj01tdVzEO3BDQMHYDjULeqpWZEQq2PH/V28GecElqKIUIyrGKdi3avZMSITBjO8WLWX6f2m
jzRY69+58qldbSNl3YSXN3n2l1oFEdIwIP86srqffMptOjlv0eIKe230XxB5IUcWyNnbPvtPo9k/
2DT64/46DhrC6ylWTiBeG/EbFhh4I5GIEbI1jg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45600)
`protect data_block
bs2e6RoThweoz9Go5JCr+QH3Tpvmtg5mdGWSsMBnVgTi8cho65HXCGU1MZ68ACje0QeRtgikJz7A
unloz1jx+N4g8RbuEf9cumCUk7gGB8bh/eBd4zppLx3IPmKrpmwtDC16/AASk72mycyQ6OFfqK3S
BpPKzs09HzSr8iicmh2avsS6JvgLWynvRS3JeHg1fTUV21xkPML5VMsRszjcztZdiFHSxvdt1YLV
SnW9pU/pHPAhz187tNTcGOh6ds8O3zCxtPH2oPoEEAf0Rvq8EBbnhccZ4Q1qqTLHVpmAGA/+pvtl
8kB8z/H0IXFt1287mSFX3VUo6GHiDBIa8qanZepdScmQ4nrrA9HWi5n1+gTjt7m9cfeuu1w3pJow
GEMFxBQmyTFrwbKxJk2gjzMrV4HkwdpT1LhhZOdB1gmabaGX0/u9jOmW+meq0ggL2xYWVG9h9+2D
CoFWDuyTqdv8SXjgakHmXgjfH9tW/+aX9g1kp5emCWBe3DfZFccqNTZebG9PkkWu3/0g1nORZ5le
FE5IoJHihzsXzXvZTsL2o8W6sXVgwe/Ct1LlRmLklibfr+YRhDkO7BhzC74Kniz3x8xjLrYTzDQ7
GAlwZxkh7lR9TbDWUdLgxGdV3QiEZbAw/UCiMgSqvJKNP4U531p69/aFC3terT06HcIBfk9C3Nqi
ghX4dYjxZeLaVyL48nhoPOc5SmIDUR8R2uxhDURJyjjvUlvV484A2CMPaUepzWl3FZMb3zU9CbpZ
/ID01u16LbF+MWU8USRhxo0ikec0r9TsTyXSoazO1ZDrGq0yJZSFIifvL1Tm4mRXpOTnh8ZiSNNt
D9lLUUJgST5809JkboAiIw/9JgFlkit41OHpLGi6+pPeXBOsVwhoRBrclb+3iMdW0xyLAsc4XSqo
EgzCTeSFqt6y7ayvSV+rSue7NwJnJj765n50gkE40hfDyEfP0OVvH8t0E+btJPHuUfeSiEJfK7Om
AhN0Zdgoo2bjnNce54xFPBQuInD4mXMGM8ttXxCMgSMuBhD5iDPq/AFUtyqVSVtDbpEMi5eO3rX0
jw9A4xe0P686rp/M5WBdwm1lHOmn0/2RuMKHPffXHq+pH2nePIcUKQMrsbgl2/4UyD20Nh5+4Fxv
7j/g9rfCiWTZ3jZdAQoTW9SVSxupMadyDG+5bGnWJeNSQOS60BYa32SLQhVI5BhubqfPOxkAIIca
ZPyh0CCjEK+razCtuZeMc4Dd9IgkQpKINaZEFGqaVLwVvTwyEMXYVDbG4dCbVGF3VJd78pgelIwQ
+IqgBzs/eFzqyx+kLD6Yk3qc1iCKaIKXQAx3eKit3FChEsgFS9/bkc7jq+WdUI/kn0kWHYinFmkC
GztFhK4uB5yj/i9v+uamtABwtjNEherxSbZsAteVC7OT1ljjbwU3bJuxRjnOe5aGwhuE8yU8Xii4
5S3OgTiv3T8wdPmqTbzmZas4tJhSlUPIheHq8WjARiIAyD0NGTsVzwlNjs1oaa3UAyXtQpHJ9FJP
fwlHCdMBvT1uKZzVS/9jDuIJzc7cFa03kyBJwQBIbVg7SZ4LnzbJikYHIzJDebt8NBnKashBPAoG
ePgWgyu9xfY5ikCbcaoD7EizNRaWXHz3jPPXduRirSqa63C5/ujRUEBg/ZBbdb2o7ROGA+2MLyM0
ZPbDbndpKRZnffCzbQcNKXWj0JZAILlYQIMX5n9M3We3isSP3+OarBIqIYt3+9TQhbmtBAfOi3a/
N3cqWz/1i8dfxBUCM8Is55xndHRJMOWLxHhMNca3Cl+PYl98Zbc24jB7Rka4njsO4ofVdb42NdBl
36clSbV1UQrMLb6lFpgJgPEo9F33p9MXoqLjx7GGHYRiVk8qfM4MFMXr0L6Varzw3Kn+Ndun/jTJ
D/sobjf/G1rX6WHxcI8/p91liPPsNPUqTy5eSpHjXUG8i1jVaJGFOKxKF/9WCxecI3ZxiEJ+mk/f
Opmb84R04+g1LQQ0nhC3BejZIUIAuzXJTJi6f0WSuQrsOADJfXufr2afFkgDz3A9jS7vXUCDbRZm
XJ7eW7JB0hDgZGZ1oaEvuz3vQymIr6q/9dhQJynBjEm5LW4xlNQDtkzkpnGzsD5yIjg2SB4hYSrc
h0MBXaRquW2InST6HNcd/N9GbcXl85YYHhn/Xm/URS/Zy5BcPCSOtIGhyFtVr0kxSYvagVgLqelb
Jk4hOUL+Kryy3oZS5OUZXycAZIlTH1U7HrJ0EjxzQI+SXnDenvHg3dPjvSxPPzozxumsDq3q91JH
8S2n0iwXkS7/wQTEmtWnBuO9pN5UcYtiql0wzSaRGf2lTnb7zjfAttWC3b+WUUbiXvCdzKjOuxyf
yLz6mGK9hVpgQUgog3ej6qFmZ4uHzAUFxNQk7JnGe8VD7thDVvZPrUJ2izzIzzBLTQ07ZldiGPHJ
PVkKXN8YWFDHnlH0OB2An4dZJipOHvp4hI7e1vRLjKle/p9vVoB0QGIo41L5+FGFaeXMdL5ORZhY
/0xOUW4IonogyWcVnzoduZjIkgXjd8Ql8WnJO+L1T4yFD/IljM7QzGt4Z1YiaIA9bTc+SnYFYG6v
s1Tz4cXRkHaaW7NxIEoYlUgzJIsFQpGHG9BSmCA9GwdC2xtWEA2XpHBvrIGPMw4rVDk2IvvXSqPN
j52fRe9iRqlwQpXfIfRtTlb1hCI8kMO51gptvN7qAHj6TFIupIeS2SEg37gBSFO5Mbsv29ox5A9y
RAYke0Znu0oHoPqohANv4i/Bt1WlfCslbFZwyDqdRXf+P+aicwU2SFtE4JFDcPn1Ji4U/jXt5/9J
7o8iCpgEwu+fRWaM5Z1+e8JaH7x3HqLo2achTGt1la+ptxgKYenTqJ9+Dlb6D0WhMqTMsEmNilPR
j8kuJul5JTSPM2U96NB2egVpg0M70q+xuWjuO8xffoXY3M5F7GLUx37jSVoD9PdtmxMGj2tuO30c
NgiVZj8WNzLhtcEAFrVf+/1BOnsMZWDz2aDQiDccRKUMkq70bW+9XsStWS8EBRR6fwf6F+e7jPY0
22D9Y0oNxOjCPeL6HcMpBno0pxIGaztoT3uhWfqJ9tznQ9a7sOhqCmayNOoxlQYVuVVGsA3r4DTb
etbmv6OhcVnRaJX9JRsYmOQeaYDACmB3giiTM+QxH9IxU+fIMD3wfNGuxEECZaImjgiZP6gUYo0I
mK3Rf4gqqgJsjfNidNVLR1/hsQWkJeQQWnW1G2scaMZn7k5bpWHncr7lfGAnKX9WSpTOUFfPhl8b
E1NXb4sgpneNX9XyE5I9H1klYJE3a/vxoIyDC2xTb9vFWAzLPk6QBF5kpUFP0uN3WBFjte+zfTVV
EhzheP5HQOneU7AKxy4eCwuezAI0/TnuQu6ITfiYO4HmpNnSMchk2g8U4xU9yppS2T+81NiHbwfQ
mSOmgtkYJBjROwwPIvXsuOrUAQrJwj/hwsDu9JoLbxi+RbeF7+y/kKBa3lj6V4GgHNmcbHOkN5oJ
wGqYCBdxqd1SGYj6trIzGaoXt5fZ7RrigVPoiacsBaJX72QDPKNMF0oNaMu5lww1oli5Givj7H66
Nzqw7O4gI16utDbxRmDvcA/45B3Bapk/EYf/5T5tBhIKy7ARBm+TYDlGEocCUl5HRVes2mp5JNhK
sARiOwJghFQr5ApZnmqiQx+FCc0+JRH8wEA9CBP0wbK3Vhq1C+wk7KvccHjLlun3ugA9lHX+QpDu
G0btJYTYUoTDVCS7rNhzzFavwmUhiX940tunLUw0c2pvWyDsOtEUd3rdTtf802gTK9Hssyx2bkli
wVCfuwaXODxfWvWMPpoZk9Chn1jujY4zCwzT8QRNr9/VfR6nVKUSMapODBMd+snrIsPrXdT5dv4n
bHzhO+VHnQWkkZ/DpEBU0ttxADMyuiAV+AGnlqK1K3ORDWpX+DH6CbYM+2d9lSFxAL8cBUMAkYsc
CtII5KiVDdeNwRTL7PaMJmdk98ylJjpBkHDzgPKlVQVOV3uWWs+Uy0fWQ7NvtQwf+vMiW9F1Ofhb
yAY8f5Zmo3IczXCn6akZIGH0qT54LWImZl42rA96KHr5m9Le/HFBrg/vTyFvaLtfSLkx4Z09PfhF
aj1LzpMkuDgDuCJfIuCLMRNtJpsuxcmFQonP6qTFd7XRX/EvmBGcRKNxKYR8CXts65hT0bb1mRrZ
2zw/pIIp6IO6rzfoJHwH8PdUYW73tQ0NQ28u/BATLKJdnIXn47jDB9ACbwoijHck5SfqNNwbgNTQ
gUDUSQItqqqQSSwwgb8AxGeqOdQ1vyyY0HDpYzYWYKFuiDmVJGBuhHe5J1mgfSof4N5vrw+nTopG
kBlw/dI8V1o6u5cQe1Upq5Lc9vr91IYY6zaQKPYbPPt7XSfLBWMAtqyI58uOCRg+5x9pMmJC1GEq
rUJ/5DJ1T1akhkBf2/VA8d7xFK4hK+HpBILISe5USWIQ7eBsD2JpH8StkRxaWYp8B77990QqMoJo
WCcb2ey+Pb1mnbMRWSzlg4Nld0iWoRPJHgJRxZ+OMxd+FR69n9PpL/FfRVXWErE/0NkCEq5NjyGS
4h2SEzE0xnxhW5pW8Btnac+Q8skrTcRYO1dw4FQ0fQKmCDmU4yA0k1bqadhG7892WcHim+itOn/4
+iW14uL3nc0CMJ13qtZY+TnmWvhy1QUP4w+6Nn8adr1iDnrd1ekCuncaAra5rxr1ENWI6A+nOkEa
/jnj6vs8PqSRvJ0w63vLMDjqfdIWG2MddGvTPXh5G/1XFICBsVEDJZvB9cwgpXvlg2BGnwYa64a0
az9BBB+s/xH6Bn/cmuTAYU88ug1UHkXeCjiNu9YTDsFRGz3l071dmprxaaCzEVBeUeLbtdS5R6Iq
NOySyhY0D5l+Zvg3xyuHEe9dDlFpHgvILAF4eA18d3fp8sP1a0T2IqCYA2JvkrHzWc+hedqR8jYD
qgQ/fBO0j3TZZtM/nd8sjRDOXQNJPSxcN/KALxMmt3nZ3Qjziv3ygb0j3hmv46tgrFZN/zWPcUkg
X2htutgUU/46IaH+0fJk0LB8MSMQS74iOTYEsnd/XisD2bCQcYVxKUajrtScxgPx1/PoTAHz5CMm
eV+/do0Xf+UXmzdtdD9Ginjkqh+NTTzU1Za+py+L81au++vHNRtxHg9MPk4YQ/sv8aMXdjziAVQj
QdXe7IKmqthiDKamv+nXrnuXr+kqOmE5/UMWM3xC1e/EGQmGWkqEEv0gKqJdZdkwi/JxepdF9Tuq
tRhRu469tgl5zjg3N+P8xHu92ZUTeLKMiH90e/pKDUQT0MP21JSgC7ulr1Nvbdw1eMFVE13zqzoq
VzOvAql7GNY+cfbYkPLvzXu5zNO/g92j2XYq1zmKLcJFLnX57wyhEX4Ag65eeujCmTC05OpHsZQO
SbmzofDkgilF0nIuarvZHongZMWT5wJOYOCk9kG5XuwwZnwlU4tWIH5EDgg+3Su93MAerw70HVWI
dYumSH1DVXn0grHvxIfH7W+I9oOyONsTO0qu+0BszCAUTvO0KSkZ6Wr238nvB4teKL40aa6G460C
Gd6IQDohymWnPstvBvIhOvwvKu++VZFvxjeXCxOdrmNrHRr3ubvTipm7k7A5kwtCDvmP/rkyd8Ix
qo6KqzDM9f3gK+jsPQjrF7lGkWjLmopwZxGl9j/ZmCWgTDl2trs5DMfeRiwveJ/CI5bwn3oVRMz5
vhJFJ9czAJiA90mphl3WDroKLjl4zmTmm90fJzsncmcztd7r9WGFBdfdQAmrRAAqM8vfR+LONgTU
xgFSegcrgq5r2Hvyzc8zQz1/vUss1DcKE8Rxagn/aPpgataOGeT8sBbLD6toIUGW3KQh7ZJ+jfIl
ke0Iy/AM3lmV/AXeRHyErOixJpKJNrjNE9FXHmBH7+gXI4n729eq93fRCbI2XQaRgk+RYc0WOesk
7XG2N+hX//NPe0uvAXzfFd1PnwLeucKVMEbmFVJ63Oww+NgkEG7ufgTEeehPPKkirVtX10bGpH/R
euPlNVVOtqqniY2W5XS9EJCR9q5aaSk/pIl649nERzw/zPotBafgTbEsCxr33GoTxs0zw0eTTDVY
ARyHHsejDrK4jKXHAjGwjDsSg2xmTVKM/hab6CUo4qI6fSYE8q9oWaxNFzI+ovMQRdz+fvO0aK2L
tFEVoiasCjHootrM/zRvh3T1qfD3hqaAUp4/fHK6LbJwhBllrtIpdDByZC4NibhnksnSQSu+XCIF
w5ivHF/zNI/um9kdrfXZavG/KuBIKNitlcvE3cYwU1ftE7vVTirdcvQl4rr58umkvLNm9kDZTOrj
DUopsZXkbSREF14pmk7QnVfL6lj3b1GG+5zbBxv3jtPzcQZQ+CSAkTm5jiIrdulAnplSDnjrLNRl
X0ajlkebArPSCcm4mEVKtTbNien3qBrNu1qvsp2qBgAvhVPe7poCvB6yCEjHLOmyW0xoZonWWIRX
89Ch1vdWP3bbGqDfpClg8PE54bIZmFklNVJKoHCVvV3L5ugHC1oNVa+FUgF/XV9qNrw+YaTJAKgv
DeDIYAIGUD+Rp1SO9scyHyYCob64hO1fGJrnsWfVl0S+yXFwtc9/YrvY8d4FcVH1FmzsHACaJkRO
tbuGiiYK35rTZqfZzFjUjaoo8vVN3Z2aUFm6nfZ/qZrZ7UrSTWzVLmtUgDIbm9QhxpDsUOzRmMKF
xK9+ZrveUu2RDIhmO64M1/9dsyA4erRNIdfJwo1mWUU5+xgAhFGtmlSxlleAtqdbV3V4jlQlsdUU
HzpbEiIYEHOSG+ocQ93bcOp+gvmsOcJq1JZjNyaiqNtxGf5Ucw9nyKJyPFlVJxXAOL0KNXZaWqye
vlRNmxWkKzEBvitnc0tUAPn0fEl9kyPr9jw9aCoOpoQqTR+YmiRJBx5Aa+aqv9izsO3UkUW6jYwh
936YKNarP5Ttg5smM1uMck3r+XoMh3N6Xpw7palRhmqr0iLCM4QN08xrrEJ1C7Pg71KuK0BV++x6
Gfjfaq8KrzwypOkYefOjK/Y5LvOi4N33mmV+bT3/FXfhL8/1dxRALw/1zbnQ+5A/cjoM4j4XmsZL
WCfG+LFACh4FC26ebYdTOboGk2VySw112BzJ/sLvWKxcGNsibK+NW199fA1Ru8OPY51Za9s88uUC
Us4ONj9ToNaHQ7ogwcw9bysZezG90H6ZQeww2OTdNEG/EUglY+pWRa58j79UWtb2lunqJgryg0SP
8fDAGGSgSUIRQb2RnWXZQ1WVKOBmPiZ1nlLbDzNdVM72ERCQCHl+3R3qeECCQ4r9HehAp0kDenDp
7fWUyI+BnOhHTP0RN8X4JApVlnIS6ri+2eTVySwnw7GBIFhgfnFNgN4Xdae0fF4The3sQqs7hMNJ
ZDv1rPY2PizJ52iPl0ruvHCgO7eclZhvz5HmEqeTjRWS6+0aFmZNMFVtrt2hO/vKO9BY/di+cjIR
9geqMRKl8BRDedRhH7IMVuw3EYV5UUCsLTEZKeCsA+ldaf7hv3q/WHlgODYoNmtCZUbw6WFhOgCo
5Z5MBjPlRI4d/VeQwAgBjQfKFzNVY5EBfQNxSFWLjR94jtOifgoCIKWvWsjVOY1cgsWdia9MqdVY
RtpMgXAgJTDdHgeTUScdqeKLzkqVLif19ZRdibr0EMzT5E22vtzqjD3pm7JMvHZrnKf8AytDLLLt
TlD7vHMRQ1zE9AEBf0OuDlNy2DLcwfvEJ/1YkbMoBfqRX/7EtBcnm0j4d+7wd10Klegu59UCgOdS
h3Ki1XgbckA6YlMBT4X069V9EqGaC+opmj8WvCFz4hUe3N84iI4R3p5Eko5hTXHv0ek/7Sw25K/z
CbGhm+yP+YHvmaHqXDm6fitQbeOrtBxVJIE2mJ+5tsTaStIrpgRqhVfOt/HlHQ/2tazhx0N4Uvn0
j6u+kL76Gz9O/ppOoaVnUDlq3Wp+2hSh5ryGpa45eh7H5+UN+E/tnLPX6eCeJfm1AsA+sxnUJCZr
9jD6n7BG1y8Os/EXKBnde1tEbJHojEi1L/ut3IZ8cV0AisaUXtt1Nukobyu7acfbcY+9Ae3ZY9oj
/gXwpCnyPWUCGSeLYiH/XlOO/EeJkjeIgadGSlJKk9t/E5XTXANVYhBZOP7yWqQWexX9Ru4W0KNo
aR47/micu803yY2Q3HfwGRZ3eWPPLciyJJvAvQxcLuI+onFcU0y/v58XBLvG/q8baL+ufNUB2/wb
9So9mMSrQvEyvNa/3SiCXCthHokw0Qx8iRlqZCIkAi4oLdivpoQYAubTDGDwLH+2JzzKUL4PiaZz
COxueWpmbc8Sehf6JHNAU5CzxjY0UJSmM47DJq6M0DuWeG9htx8wRBNwogzpZmFWL02hikB/VDCo
1EYZZWKKSot9iM2dZ4djgpor31kGj076ykFuZCyyeuW7TffOIgARLX5dl4+gjEc8+Sfw2gklsJ68
LqBx/6s9fKyXOVNU9TJzbz+sZ8YmYK0IZq/lxX8VIJixwt/3YxoMqVHndlM/5/LhUKWgsO/cPs2Y
qYqpcwuQ6EkbQo/ikQO4ZY5sx54m12ZrDY4ZP0yMcPrd+HLtQcjAXRaLPuCN0c8YlpEjCIyY90A8
85NYx6qPnf/YL1pQIccG1p5YJ95fXfryKoHixQjpycRswLzXbXxfHudMkBYjqHOwmrgrSpRvAbHZ
dJArp6aShO7XkVc1f+6oX5EkkC+tJ28DDsmW6ye/bLZ5jBbEsbCYSkC7ui0YYxhrFkBxyFhdNK2+
S02JRUYhutHyS4QVhBj4Lsq7DH0Bt8vVj6U1x3c3QBgPSLDxcK0fwWkpjvLPtldxqcy4sgpog/rO
oIbdlm9r2qHksgNRj30HfzudiiP+yeF8sJQPsS7vZieaBFy96+bhKyMwHfaU9mmr79kV+2tg4AZA
LWjSwCpIk0cZaKfc+8RdNaFRgPVu9h4uUWKfYebwfLE3sW6LQFRS4f679vlTUgcErvYK4/5AyZWY
KOiQIi39ZVrTaUZfCLpuSB5cJvAj6aAD18Ffgbww7euwxT4SpsCm58rZUeO2cxKUBD/f08lBW0ms
SSHWrRBeNpOgJk+hMYPiU9JVub7st+YHDr1Wwi5iAU6csF4/0t6fI7aU96K4EMVG16IO16Ju37av
MPPZuhdLly+ZEDBLQPdhHeChnKxB14D/GEskHmNUCooaiPadu+MoFiZZj0F8HXNcC02znBs/WrhH
wseBHEPE16J6YKiBSPt5fq51RkyBhfdZ4+Oz6jWUqGce/h1/8kvEyoC6hLPh36zrpJALxh+I1zFy
ENLdc+R8G1iAmkgTnrcKD9ybaHCrAHd86zlKGFJ5u674cwjqVD0x6wRiGXYU8UrwLXbXjqxF4L5U
Ssu5L8h9mKjLLQvx3VTKn8uU4RMh7SxKXP/AjRJmqUPO6I5zDp7LCrPk1xqYriE+gaYOkAcE7aAp
/GTpMyZ9otybbM6mGOzs9XZ2C2YEGfS4Wwez1+g0T5WBCj/icgcG+//kkiH7UmIWc1lSJ5pZRcwX
7WqIrhTka/GGhew7ycDPQ+gCrViFPBXhk+d+8ohhrYBIhQ00rMqjTfmJy6WtNzqTABHrKfBJ9hVg
FWU2xHJeJ7XqvhMtx7V8vFnbvlyC3Fsytahk98Lv+oCrg3+9oXVp/e/vLjHNopfFXW7qAYmY1YFd
X5mW8MWbB0TE4huqSt01kPAgYdrqwkvUCsMCjVxI/Ea02Q9xxGdcHR/xsgpdSOzkGoNI8P/bUPO5
QtHew6iuJx4aToZh7AKSPPGa+fQTlzWOtaQhc35smiVq6nNpleI+g5iYzMd/QEAT/SdAosfryykw
Yt3xVsEoFh08/59TrCj+XNzKincETFKV5/g7LO80YB6nh0N3Yjj9UK/iTdlHr0Tf4ReSSa2NARIU
jIB1VWxHdINhZsCaAdfpoVL7UD/vOLU+PUUApVK/5cHPTMv0YJ4xTqFiFxj8IxAUX9vN+pVy5ATX
Z9WGFL6vMXX9Zx+Ml8Bz8I6JynOzLG+5suoT4EgYhV60l5nvQJmPlKTmPpRK4BM3tWgeo+nFEBm8
qZxXtfnX4eNAhhWjK2cbdrHz3vorvl3alIHBohbeKRSrnNx4hBNsk6mLPGkBxl+lGoLE3ExM0Der
I0qqfwJp+rXvs0fJvmR67KU50+5KEhADshRhQVtRtJ+tmyZaKyYz5LNUWJPq2Rp9u03tmt+PqLGx
QEJIoM/4wWKErWYYmEE1hnhSO51jT014nFPfv2I9FY4FXn7NM/jV1W1M5KLHwKVosT0Zdg/IJpWm
ALZ7zA0/14GeFCTULV6u+J8lODsrVzhxgHCPv+JRuYu/OrxdY0KoTQISqxrLnd0vsvWmSe4mNdyZ
WRPCer0fDPJHvGe4JRYw7ica2shUjvIAx1WDxQNHZhCi1muUjmUSfCFW40AGW1KWQh3N5DYHczCq
4dS9CPEJ/2HRKtnL9FhwHv6kr4tRx76/1D5VnST3Y6XBBqYsmI258+6OYDgy3Da3OEoUs9kiscgx
9GOKDaRzSQMF6Fk8tJhaj9YGzX7HN1UKCMV9xBhlCIz37H4fC/h9QMgnSizxYFOvaPwh5SKsYXp/
oQ5DC5++IvFKLA1Dm6ZABAPVwz/qF3LIgI5tIiYhVxMMoTC5DaVRm3mfuGZX24nRxKdnKiVoWyUB
f+vftwHAOAoMAc/gL9yuXKPHQ2VU4JMwgMHQLw9YtgLxDjpoldBjrvz2DC185Z++7ISRDCt+hTYg
CyaVgqJojI3qaUI8+AdnHDgAR27FHq0PVkAk6PHav45JIwV26Vv1MaD+bgRCdJ157ZW3HY9Oy/3H
O3YyjKWylTFgy8lVDTtuZsU72S4886mcBr7porEJMw2JoYqgN/wOQbiFy+SmqO73R7pWpAa65Kea
oFd9QjoM8r5KxZdmH/KHHVjNTgmX4aINgUq7VXh6YH7M2A7MYQPuTpNrp5eVo2eBr4WzmKGFQnuD
RzsuRO+1M4h7N2q+gwVPYiqSkDkbqwdL7RDnl/8xdk642sAWY8lvqzFfTrtjoI7aIdvZpZaxZi3L
tGT+FwvUZ+MQxlqu7/51Vqn8cdJ6/F8cGB1C88XjY30KOG+fbufBa5jGINdlaoSPdy3QR64DXAo8
WoYbmaACDsCoR7apcIY3belT0d/lPZ6aASqrgxmejuLfWZP7Cqlsz3Hsu4Ha5Uy3RO23YhP79SkZ
+XB9Xn1Km1kt7zoOQZ/AqMsUeiYR9Ex/23tjiJW9oIPIQ4EwDypWcZPAdfXMTuz3pfRg8NXiL85p
1i9Iw2AS9OoluVSKkuqeUPIt92C6Z6HSdm8JnXweLKu8qyh/A1g1x6G5Yn01GztttowvEDAnAFu3
3ww4W3Rg19ij/UubjT/nlfQCHdabqShX2n2PuuL/8ryr0WDo5xr0sJ2fiJwMTDDGx5KspZX8DMbt
hxZ8Bxz6VdbVEXRV5PGGSCPcj5p/L6fkIHZksPx+sHsSIth1P2gRZxvItGkMdT/4TpyLRae0KXNL
9gSzXVEABLyHCkvU5K12ha8Qqehi4wWYiByllsnyLM0SyPMDEPVOzEIJzxC2NSabxNcucf0oeG6R
P6o7+wfxA35+vW3J53GMnYSJDpsKaT7poXrVObY2cNJi206vGlJBrTCDogxMMvWtcxbQoZ3MCwlL
GbeItOoQ6Cki5XVWxR4dJQjdGHgpssTPUQLp/JOy/36MT/BqxmmL5AzDov+g5AoXwiGyCzUu4Kuj
9htBTsN76Fl2bEETpyGhzhbUxlbwAhYhrfiSut9fMyYxb3TLsX7i7ZNBc5FNZxC+5Mz4lepiNceg
Y4lPP6BtIi0tmpw6qydrFqCAIfqy6na3ZS8JJKTI8rVsffohm4y7yWd71aNgUDa5b9JXwiOWHaJl
JMCvccMVlxWYCL6lRDfPZywGfmzkB3ET7+CTurSx7/a2cPCT/FM1DMcMruDyxt+/47XP7+2fduLC
yBU1fh+UkeIuQQOruJTm4JtrVSba45cepMWtc5E86sRZu+qUy+rUauqkNC9cQ2U22yrN4xubeJPe
98fjEnAWSfMHGWd9Ja5KpJtWXSVws0HEJ+q3NJuxVeu6C+vLwFQTtAG3b2pvrs1q4c5hNMNpiM3l
zq8pJT5Yjf4NNR6AN9P2ACCS4SJ7MvnBot+2DqN2otWxh5KizQnoOhliFecVexd5ewGZBlaPd5KG
M5VqGXTnj2vBB6Y/F8nQ/8gk5b5QZBnUycMoKny4my/MTApyIgI1Xa8QFyMpzv8hqhRWuVQ1L0hM
8+BGLoatWxmCbuRFq/QqCSjDJL2oT28Flfvantfmc37f65Z6p6SkuS84gXFxes3db3/hCnS4MmGa
1cuZPJIKfvw+RPlRAQVrhSbVaZHLZlR68nqdm453k6EHVOmZWzF1zWHpqJ7ETkMZwZLK+Rml1NqY
bnT973IQdOqYhReeYN3u4MflkZOhkbayZ8WCt1GpRN/tyg5nCwTnuk8dJLC4k2zNpPBFzLB8d2ZW
WoaDByRMlIRGrloc9nh9/v1wUgO9IR4mR31vAsS29LUtqqi8do1IXqyi6YBNO5+OPogRpa6UFtdS
YLZ9wbeY0zjHewhC3u0FpoMqmfz1L4Tr/p1w3C7p+WPWoyrm2/fcCNWOMGAFKPhLmLbejIirOJDX
t2loBbVvlU2+6h/f+hL1S+nT5y4R+CM5YROOpm2jsp7/h46377uD0J68L6bCJ15gYnaIp5L+kZdd
fw1F95uQr5SA9ovXxdvCpZcEMrQeJGVMYX2D2bG6vy9Udc8gQh0wtdChqLjZ3hXzAEvT4JOXWW6I
ayLtDn5AIuHv1c6ZSJM/buxg7jHqq78AxLyfQFD+FpkfNWAdB8mme00Wf/xLT/X/IG+yinm1pHVv
ZR6QQ4O7+PjTWW0/XRkA5SGm5eHmXVI1H8KSqS6KOM4waMvqNqaa7BIS6SSD240E86yXEl19hivR
Zgc62iz5f81Pv55/nJMFbfFFrfX7cLqVkCHC+/q9+qfA75wG5G4zp3gKI0mxCuy+hEk1dE9nTZzj
d0rqeP004GCSTfwxWgWWVCI/jVDo1Xb8RmmLsEitZP+CvyM4LYuqdOAL94HKobpSC+4RL2SYwAlx
9z1ZPVB/bFl2yAy1QPMQVPYVr/9BLEvnYib49IHry2pXrNEMOhhXvtDqnMjor03tSSiPLdVsjbMZ
KetkckS3hfMCWd6hlznQ0FzKGZQQw0d3Jy/igZ9GsoSBkk2lZYzJ8CSsM7n9UOCIZ85KgEhI9n1N
oci8S/ps3/Q943r5Xf86vViQOSw3EnXzxb9vu/nznU4zVoC9upJAnEx6Jpz7HcJSmun9uNRyMkVp
KurXILSwYlOwIssucTK5l6PKwAut21a50M7VBnCIHNOvGH4tZSU+UnlYrkoHY3iSfqe334tHWmli
WcYVyz4agWKmFkC1si+HpbBxBNzCvst6Em+5kr0ngyk5je1mUyOEdJccJ7iQAt4KiKqUaMvIxrJO
lFhU2l+wAY/G6BNeTb6EKARsgzkbEk8N8LRIT5gYVYEMet2Wjk8tz2Mc8/yT6NF55CtouVamS3Ws
J+IPGa7oIf/5UDSdNw72I0n/QtEem37Mf1sR51oZYwDjl3Y86XN5IP5Uy91I3oTnkXOBmmOWSXnr
GZgnUDeQKNmx/arnMg9QpEfn3WoEeo4SIu0Neav3kcHsmgnYjoge+tV/9nkAaIDNwQgkOQ6u0u6/
cRPGetqaf2mWaFlmKXezRbjq95A3+RTHC5jEl5Uh2q+haAAyY4nbHnSt9EWPk/gEDb+pBtZ0Wi4l
NXot0XuqRpxIw5N1gKQWbXo8b8ScVaFhoC7VoFaUy8R2zzIYl40bnQbzNCxCv2+UbdpG4zwis9fG
vao7DFOMDoBxsFfmnq41nwjO0kU4tgChykMoA4GbFTHMN894PrTrHPCdFqeftiSFIyyWFArAJwn5
ToWtqqvctf5iEQ5LBEnyUtz6xTgU/IuLAm8t1lphc3mO3U9ziLRnwET0vicznBBOqsbv+eZGpieS
NZyGrAPb5T3xp6qWGl0M16MXO4o8w2MUA0hcToZjniUhkx/wtNqK/mDOfPvkmHC8fDJRYP/jMYdY
Sv9Xipz7KjlhZiPvOa+yqDa7ZLHg3BpdJzsiQMNFFbaYpKv/RlCXFkj0sfQniLqZJgD8enGRsIJj
eUXGtkAxWXm/awMN3D4yF6aV+mXAXAL9TG+043Mg5MhMKdVG8ahoxWy9eZIoU/BKwHaCP/dlWQ73
usxa9TEkZ+NIL6S2n8ECU8laH0a6MyvRZnvGG4mqGTHs15lI20eBiVgr/H8XURk6QF2DG18KQaFc
rnVKCfXgs76bbvJ1NBWIsiAg9stZHqp9NJYxoKbKtunM4JV21c++d1bs20M4wimJPnvjrtmnOaAj
4XsDsbnbNFAEOGXarZEve20eLVPGv0m6rNIh1ukMJesZ2WoQrZ/XPcVBppAapHZjW0DBTy2B3jme
16YWhSYpb/58ndehjaaoHh5xQ2EYLjwNEY3Zu4a1ikzHcBb7l4zXxy1XKMqg6dKUc/akw1Dydypq
ltZ4CVAvN6eTY4g0UuurWkb9KNQe79FSIV1c15XMR/Yny9j7wOv550Rklt78l1OLxPLyUyyfM260
vAaectC4IpwAFdbJltkdHSu8S3m0oBUoZ2CDAz/hTkvQkgZuJYtX4EsTf1rWbTU6d7JWWZcYAvSR
fNlgzNzgNHrZzpynQhHjwhHXG6oJn3q2tLWZ9tjeBv7KOQN+1bNw/6dhz/OR/UiW4eE7YfORR5p/
DXd9oBfaxZwsc6a0+5q92LKNC7DgMx1Kz8wHuu0TUxPablwbVXDwdlyJJaSqpqaWfbbjkyDgNRls
cm9JB2uOBck0hb9gf/hPckhsHjKl1PlAPtu/X8y/i2eZZs513GldMGa/gq67TkPNNJTqnZwCVSoA
qwJXRxBVOEB2P1DA4ex6+PM2CP9nL2mY3NfabWotbt2PByg0JK7//xg1mPvrGNl/wgWZfB+QAsQY
qykuekHR2q61zepcUTsMDv8kae82wNrSxnHTIoy4O0uutVVOoSgt5nLm5qbeQcBPBKhpp3ZZscT+
C9k4gojvPWPF1bJXEOdwjn95QmQqmxYqm/Qy+L+yPOYSVMPSqBgF0GnixuD4tB2zRNt/UJf3Sre+
URhzK/qlbA1LDLQQhqwD2R4pYjcI2/wj6l5SvLJ57IQkNPV7ABcFDIk2ySPiSObTDxe3WiXejv6M
t0BUMrueju6mKD2sDcxc4u/O11SybCD4ZhL5CFsV4FvjrXcfOnUNq1rqwF30sldowoEkk63LS8Mj
F7Kha7wB0MAabGAL9HjbN35UJ3RDIlE3Mm2uokewe+jJU8rLR24GRFD1TJo50ieRXa1lvw3qtN2z
kHqt2j6mvTbIa4WGriiia5l2kcd3dW1521W3aGHS+zKXz1gRFi4vj7jr9mRmzpCz6GfJAKuzSMl0
EtQLHxhrl3Uy3+RCxK28KQ4+l0iOQafNg94eGFP0KHvWqZ0OPBrB7rTdycv+IQ8Bsaqg9+3oJTDu
dzYVPrRoBMnO5CS7Yo7zV3z+UOB3oGpygSBj6c0FBYbpmJp5kVcFteDztv+t9oha24Q0Nw02hfZb
CLBD+axQ0jgurCfCBnB5d4pfLrGeBBrdNRMqfcqMKLb+wx8PM4+VNLVyWs0hnC/C2g/5OEVDheiR
IA1XWJggdyfeJ7TAdCddFgah9tGbB4i5bJp1rxl7nmxXTiZjOyhQrQ50kozX0Hfhxbm7EVNudjKe
Gk9le6jY65AnSKPOlukVOVLD/K+6osE0nGkh+4LExxgA0svzHzcMGvM5lltXOTzNDtkdqb7UqoVv
bbrt3TdqcMVTH7D6THYiTiHCbS3tSImaAzK1QR8YqCPI90qke1d/qvIhKW01w1MuUuKjSmEAw3mc
9spUmMjjRDDX4lFnaXv07cz96NgCK/oWoUqcWoprR2KO1xW0GQ7u8gezqMy01KQEaEZ1991xbp5J
71Krm1QJUQNX7gt70+XssoN9DRV7GC711XIYJMQ4/jXTGP3Xv0FqEIamfo1lSkvm2vdzXxFsG6/i
1hcZIDXWS6iwCfo2iTJmT+PCBcmiLmP4Magcx/H5ID/sgHSvOYf04TDrHwjFNxrtlHuWQsiRqWBp
/QyNf1/eU2MH1LjXA6FwYZbnerwrm/1D3Mg8qEwHYanNt6qDePb1EYNObBCUW6Qb97fn7A0znxTK
9EJ3yVyO6fxAtJsFIo/qgZo06x24s8uyeNlfrJ92dI+PblthKx/5259vBOtndm6rp7hbaPGotixA
esOhz9/sicwY0d2h2Iuf0CUITet0uEjxk0SHXFPl5k9Z9HmHljLfVmH7Th6otrDhoJdKXay4TmPy
UuMCWrvV3/4Iw/KeaHRtHX9Gs5GIHQRsc+aqhiZVKo0XlBGvoMqjC+2n5EChcBURQP2FSWLcyQ3t
PxXCvSF9JPe7JvqpTj+d0OeQ3mn5kNMXGUaDlF3QoUyKr1yJRxrbGEqUh9GVssiTkhVaUfrmkdi6
xk/JYLZeoRXNj/2l4xjvGFfE+jntXBNQRlV74BGN2l4sRoE1kyrXUhqzSCMyY/AwG4FCm3yAfJas
GnXaBu1kQtIknA8R8fIU3O6Mby7kNzL6BCJAQbKCprdy/CtiYFjjgDxFsg3JihC0wcoJEm4Qmni7
wL+NgGMM7qNJrJX4s3KFUMsBlpsz5nk/eYpbMVl9vg9HqD+s46w/unKH/gzaH2u/C9QUTMHhIsW/
lKxz7/S4CSF5SRjDOj1mAplMDNTYcYfZsw52g8Fe2WlnG0oFPBpa6mgCq7NF0bnZuBzN/OsuHOAF
8uJHFIeuI7LIwKbaO62A/4JiQV6tBN6VeugHNmLwN19dgEzUW5iyJ+dxwdzCy3SIvvKG4HtTaT1I
QRSofPMJQ+7pE42Ld+zEBv98cHm3SYeiMnXbVJk5tNAzDr1V1lRiaVF3qgopM5SXWRMYhpgE5M4e
nN692qN3HHAXPvMvdbluXXa9qLnVZIrs7jsVQZew25Nvt9EsoityEN3GU3+Xu+Z5e01FNF5HFjL2
p9sNtTYLe3pagKINo4wxRBFkBuA486kfnkduRnJ5oY7gDJ7cPzxBA9oabyqrvPR5oEigNg6ZIxyl
DN93t85bJNK7IxV/JKqmgizOry7c+AIsLJ/YPnTZD1mv/jg2AIt5G6mDJiTbdwwZbXjKIc5gaqb8
91bT1r1hzH0RX75eyJNcyE4SbPXGTQVfC7TaPY8/8PZfbR6A9VZHgqOPnhLFUGyImY3o904xd+wU
eKvItmOouGSDbCC7jzqEtf9H7Wt42aMXyccuk/TLFUs6Uk2q6pHyPWpjyUW/dBryyoe/iGHDUR+D
2XGCzkkfqTpGcbv5gL5ylKCieBmxHOnPqqridmE/pQkO+/+LZxKCNajfGPhtJcKtiJWPzGOX8bBz
tTcXTuDC2lUyaM4bqt16kep116QEzam/G8ik6lLt2MvPga915PpzrOeDGArjqt5zMXB1hF22wZZT
aZw1ew9Mu0gcw4Q6wpGU2RSO8dnDsZXfFLedLdYRjrgxoiZkHblPnopW1ztnh/dAd7m4DLAdto4W
agpmm1pBHSeMx5cfaBl8um+74l/8swj08+wCHm9OZY/Dw2XV8aCeN7OayZ/3cCx2myQOp24EYjOr
rWi4783pMZ0cAsfj5XlClXOySLQ9GUOQpOlIjT3BpowisAHZ+oRohcLh55pbxOzTMaz0M7iQQ7SC
swm7ps7B38X3VMl/NoLzUKChV7Feh0aG9aSJnIyNiTwqAXE+JQA5GWFE2WHBaEaNs0r7ljsdlsxw
SVbxeh4KmQhkXGS2ZNe5eiGJaQHBymLKRcReZd4HZ+rS/kRcN90+21l+IfoRTldEq5RxHP6CxtjA
+R1JwMr4FQ02rQm7aWfoNumT5hb8x+mT6E4U3BbwBqnA/UA4yY1a6m5Wyk9ufw/g5jfRlWj8KDan
Gx42bNPZ/rVtt1LnLgu35xj5XzIpiahQOGoch02xSlDo+6b4US8m45huqwrEAdHERW7TzxwDqEad
1TMWvxYR7TRmEJYlYrbZVLJ8zbIm7an/qANI6XeM2O0YRgXB7zd13tIdKDLW7+SGrwS3Rschaft6
F/9rm69W8Mnfe6lXvUB6l5/PZFuhmqT9vyXYJvxDFSBKmPjHmQNtoSPEVPVKskG/hPKyJx50IlPN
Uni1HkSAo/slCZMKa6Xiw+AJOmsdIwkM7KSEtMU+T44HFpbR+3LuErgH1jJIN7Qau+0Y7nUK4Hfs
Opms2GjZMcYVv88toLFQJNdX4iqLzUqrqJMGfTEn4GQJJ17TY/mLIpQva6T/KNQP7bYKR7SeoZ5s
F/EISzIfcse0amuYEPj7o1Z77ddXzZR989dfDAdxSarntpRMTNHJJsmYkOvOCKF1XNVshtwC4qp1
Mk31CGyhi/hKnvh1wEMhXabyHMJnALppaWNHd64UBXJXYLYba9AULsWuKWr47TLVDARuehh7usum
0ZXDgFmqTZ/AGL4a7cDVHhXD5sLH/vR58bkVAMXPmGGWeV83geWZp8CvxGJJtTqwdL6grrBXn1KP
7F27P0Ujhp9ywOqq2K6OsoZrR/oyU7JWALuApDwLWIL7WICtJ+slL4k4t7gY624oTHziCqwkE5Iy
e8PFN54XP9Cck84FZedTXGEfN1PbaL92doDdJzgcAZC3/db/jSodAV7HWNIQ8LPCP6al1zuaauqe
ODgBRBS53JQQE7B6JQg6NwBjP4y5IETDqt9sXAU0SmelYdRpn8lQbSz1fm5zrapjjc8hWZoi6Hph
q7qemj0AHStA1VdGhrVp6MWNunBSqZuTtS6hRe9OYxXboID7C90QhLkuUZ+2Wg2biqastFUW0Jdr
Rmg/UCMtWrjkIcV1xEp2vcyCMNmmTm2mVFXtN+uffCjpxrk5kaJaTNKPyKVhrv/QAz1+5tqn4X61
rCiUgCIGyoWAdDKSDX31RlwXrbD40YsvclEOHMyguDpGFI+y24o+v29Eiq3X0HqVo0a+A/Leo8hH
G1hgXa4Jb4e+X8FgB7BfP8ig46lKTSFlwgOY7ZHdZ8TdrjgGkaugQBT400IZc8yp4r6G1M7lCzSe
cMLFr/dnQ8NC5aFOh8nzixDxcE7Kvyvy8JPsjL5aPDNprBRGVO5/hKY0FHnzvBjDbVjUpeo507r5
CVisg1/47qxMYjUwMAPUQYliBtNhT4toCa/GKfjbWF+Wo2DiJFY888DiGbOYNyxg6n5Jg6P3kbQR
3H8Lh19nSz+IJd53cZd3yrvKPgHaI8sKE6jQpsSjyvC5dR1bp17iMeFDTCOj1w7pkUMvgi/6FQ8U
8N7QQx+RJ7eG/kV2SnZ+xp+1o/Y5Na3WdbtOhnEoeTSXLOCutQs2f0EgnOnq3FYTuXljK499XrH1
zVfSEBiRL8pHDmrY/cseiJqR5CAcF37a7evb//kJ2AI/n275dSXSFKcHNOrf5zvjYRxFu/+gX2MC
vATcnggXNWyrGRlAT4v7Kd2qJK+wuK4vaKrETd4zGTd+aKpNveqrsoeTTBfPwojECw+XaV1dkxeq
6YmK2RNxCxk5e1c9rXLE72LR7yL2POIX/d4wwmEkBgOuCzxPb+dfGendGmzLOSCbT7IzhFw7Nnbs
1DvdQqp3FqvY6ScCyEL2h4GGaLbhhx8EUKiJOm8QW4wNtVD50acSS0HqOBJ4zUNQSJ8S0h9p5nzC
WxDzCL7hvOadH4bPh02TkKrqgSpg4NMKGMWyUfcmWNsuFoRC3ucZJ7lSfPA41P0Z5DDW9cyrLEEL
f8WcVyDNhV+ijJ/VN7kmFODIwS6GZuufbMNqWn2TmmKmDBtPYJmKN8x6iwv6weWpcgaaQIkjWks/
OxGDfGFMQIQooDIE3OpjvS3LDQseDow7j3uEqjj6/r6zGiB+Ef0Pftrbav/nO6tKvrRFmU1cwbLo
nPOwrGekPVhYlDBl/0o9VNW0Gd2rfJpsOSmLwaXWEYmJdn7DGsZKHSqW8vAwKTqFKlcpX5hpfPlP
YRRWfClmDi9ANpdyD4NGVv8sLc6lJ8IIqC0sFMF5+YDneJnvyByC3HtpCW2ycmHUT7V5SQloxlHB
okVR9Ya1xr8/8g8N+Dvj9QWAbObqh8SKir0L39eWuP7UWm7bq0QM6LRKOBDr6ZPuo1B9X1w2S4CC
g9KIACtXQlr+Cl3Z5SJBp8vZPIRfBqsG/SJdB5NOpTUzflSIdPN/3xD1oMHZrIFCYx1AltJBIO1O
yEjJ+GDpE/BSlNUqWX2tfG/J7tL2gvvRtRtdj4BeKskzg56Exm7QDnhx6ShnKYM9KjRh5wLcL+6m
/4V+eBJKbsNJeCkIoL4PcP948gsVvdGlrNYssnUdi7cbnH+E3QOtCUYaoMGng7eCi0xhfAYgL0E5
/WU+XHWTMj1CzIBZ3pyKYy2I4zY+BBHWC7XKYHmjezDiCZoy1gHsHcL+lVFYrXTCmgddJAwYiS8s
R1vKbZVvMo/0kKtODP9MkMhW1HkpF8heCZjVivQ6vtX9mp3HOfDUYCSVTwT8bmR72bRO4cQHmRvF
yGm5J2bDPiadRd5PKURugkPfMM2PUy8dnHzBu18YTFl3k/R3/C31yl8m/+vb2EzwQ7S+st7yXDKY
TI04Zl3TfShZDGPRF+neTWCYZzExX64aYQX0BvvjBXxTm+VaFjZn+otGvqeUHAggSY/bhRDzgGRd
jeA4n9uo4JM1nGELBMdbs4QdQ2PSHbXZmLHEMNFWKhqoIltA2RbhOBbLqCpmzmOqGIQC/5WrJrT3
o8Aw5deMm1wilT9FvbJJHKQCNJfyZuAvZwqdj+hi/1FejanzWtEnWsFAWR6RkyuTU4fT6J9de/EB
Dx0pWGHR0ROMHallDCgA/qjngHR6JNXJOHgItobCdh41XIDKziW8FiMaw4aCYQFUMdbJDRLI1T8v
MWDUlxcA3KLlPz9EDuehQszXzKmf2qMOEAyJ2R1H8Swyx1CDWeXrgqD8a1fVm60FtUntYgXV1uzM
sP8VL0EYA9ng7vnToetzO2AitIq1U8Un7sz/gnBOHeka2fURgfrU54sii93Pr1rrSKoZlwS//Zbu
sG/K9F8iIWUFsWoLS7K3CNwJas1kEzdRSJvXXJFN0FcTV00tm+Z8q5zV2veqry6iiFpxMOF+yz6z
f2TFXzcxYBoKyng8TR2C3daax7l2tny2z+uF7lz8yjBmtxRjQf/BxuVoynuBSN9wJs1mD3wVIdT/
NfwaDYA/4OhVTZTjN5whw1ivCIlxYz8E5VjDjXP+toe5oeCmknDo8A2KCOCLqzOQdPVTiqenQVwh
KKZGsZHygzq1B7oL+B1wcWMBgEo1j8LwtLdsIS7aneYkLDCqH9T6U/sza1+/KLlLFyU6oqTBd1zZ
UIP94m8u4r0KIbwLHut1aMvPsJsJgWgwK2ow56g9yl5ALu7X0wT2NOXesb1cpR5hd3+m+T73X1qX
V0KKin6WKu6A4YLyXRDFRZRIF7K/o+o0tj53eGy99/rAx8sAtMjtkTeedI1bJkzV4iIz4HtelvVT
o09ha2oIpnECCUoG/z5ztZrKZkX2FwqIDqDh3PqVNvM8ZV6OgzIAVtaRR7qOXzwA+aMxSshTCHmX
16gVfYQYMDvMcwWbxCAX0cgmYPumaCz2HT1d4FdCpVaf4ee6ImUui3u5ly/qsT0WYVETnC9h9sHg
mInTgiFNp5PitFneuKVi7RYk+AiLNFQmzRUJxiVczarjwmDO2MjWwu0ogmGRC148nEISMt5w7Cp9
day+4WFgzh3s+sAuUrGxcrxr0zfuL4tutRFukzevOtITiEu0VDp9llN2JMjnMAeUxGo7wPkCNGdJ
VC6yKJstakagu8fAHIjhp9VSsOSV3UNF0oFyPRQAlItmjzO/W/peZ3iz0SPNUAiprIN39lTzCQk+
5R9PBO/z+3cwaNDWACWnn51mmp41Zik7ML3ZLTFYo/y0qgDLTvLB7LU1VD5smpEBVziKrTHCaDv2
scPN66K9sWpG/7sHSindDKrGV5Bt6oDvwpSStrr886nDoCZw2BbS1Mi0WZaBFcPTN+l2An53Ie5b
st0QDM6JAoOSY7qotbHY6SPIDPVn8Z4YD3RvmWTfc/biCje3jzqH6GcWGos7WAD1vtTK6HXqmpKf
uQOm5nm30V/x8oX5ZOZFsJBs95GIsKpp2717WJ5IkOI/V7mLzxzL2bqKhnPksfePr+ySlKqDvVXR
+bNl4m1CDHQDtLdKnDIDwVavREcU+VkV37AvDjODkOLkylCEt7LbAL496J8TF+fZPqBHR8oFleqx
KN2193JTqs4c3PWiamsjp6ysi4K+4jqEThwZK2Y/lNmMhhzSKtv5BxzIED2jBvkhZv+atfWdhzXb
n5bhDcoOn5cpNku4+mn8OSttmfSylH7kjWEtheVM3S+9/xqimCoxtu594bIuvCOZlOtzNoC/3NbF
bI+yqnBUgSpyKY30P5xK0SFTMERhGNZ3KkZbEcOEdaCS/7OWnQn0oEXFHY/tTJkpZppN1luDhCnf
FV6V/CRxdKwpDHGIaA0Jf4jhdMPeckPjVqkbvOoI+un3bl0Ll5oSjmJoNCSvZTnH4lecI4jjUuq/
ZOeI9hZuDQn5Mx1gItjq/jwLct5gjimCFxM/n5tKtJ8Q5pzmPp7ed5H+hKRLbMVGfCf/fDkyMsLz
8n/JnhI8gcOwrSQqcnBDf6K5dpuGYYJuAGAG0pcxplLnSStS09cgRvSLJ1gYHeKDBmeP8VHpkY0I
ypiq/3QXIj85/SOrY8ZKOsCoPJprcNCZgxD90ZlR7KeMPZFtxoweKn/LfxlG4rTHLMAqffBO5YMs
+uiW1qsxJvYwYFD9MgMaH4tAOhyhqUX7Fv/5E4SqctcCChxlZrtf535RiYLlgxGaezlfc1Aw8TFS
UPqqUmeXet7qPZPzMc4HSTvpPTXVBgKinBOXjMiu2YZPvMJjbYwZxOg479SkDbZWprwSXFfyC0hR
wmWeYV+9LXL12VZQIcJzQBMj35adSzY635LQY13xVyKMnQ7rZiCjaCtCS8+R5kXorAiHcp4ecJQa
oKzevXwLn1ilOtr7qxK3D7gpQ3eRaPhFl7WyXnRPafO3CvI6E0rZk+kAYrEV9XvVOGuSv9bNWsir
0Q0lTmBnBtc3ptngsNHfZtxlQRyDX+oGpgZLIeYnyhDyRKPEnpiYZYyL/bVOkONl9rPLz+/6ydoU
1e++OjlwNlxYNhMfbZiliKjHv7RVQqsj4p0dl5ovj0wDFZtWdryTird8J+M8H+Y/cjNgSAPxYlU8
TZQq5c4E3DEgeFu1lxMj9/+nWH/PPvrI+TwwhghjFcnYs4wB4RVRaGkRgX1zzp5nrDFcl//8DEkh
MyDpnB+SdUZoVp8CCcI7/v0MoYoLyCB2lJhexNdA3bJLm0u6uaJUHAQzYD0OuEMg8nqWIiBsUlmJ
OAeAYcdr6lsGZ8qgp/OnamH2u0Rzk2+qSUqannXR4Qarri8yaPaisAooWbqqBQB/cpx2XTS3vfwm
kp7o0zKxLrnAs9u009wfPCHc7sTKdsX8hGA1V55zenFMFSig25ooReNVuDxdHRXRYOjQel0iCM7r
/mmeKUiUYDE0y4K0pVGs/Mlr1p2S+3/4iUJYzirWm0+Azatru4d2AqvkPIjALg+qntM3nkHSmw2n
2cy2u39XDXvl3MWTkeA+LDjcnyKnnsygJ9jf6TYoeENumlL703xlPRedfrfYGV5fhbeTrGZGkTXO
A4EPe31f8SRDOuRxm4ifjoUPASoKolT5SJjJ+dauCNp5/nWwz2WCLryeh9jzwyLmcGWBjk2M1gXR
4/tiAdsahnAqK4YMVt6ToyyVOTxJOcHGZFtIez23IDIt5S451YmDFV5ewJmkuNnZTco+d6sxmfbi
jF7ntVyhjN2yuFNZiOndOiI2eT+JtfiGAeD/1OZg4rQwHZoYjPCcRlcbtjmfEbv4JOobAQf7C22F
FpAz6bb4y7QnSXJrh7SsuC6395aHArnauNZ7JluDDZSkRRSQYVwptcw5Y/R2RssoS8g+WJpODLTT
mt/cAUWttxQm5C2EmLbCqfTHJBRnNiMfbJTsFisgFjkH9IFPQ+PgiF4fzHTBNut5QNEnR7SdmZcr
KsUaiOpBMHXLFcXSp4/p0HFyc6AI/7d6dw0akjy5BN9iCnarT7V1Bw7nq7zjvCHliR/KOpgtHVAV
GUxR3l8DKTGCFXsSJSfZGXa/jHrAygy5Z5eZU8+kVa9Yrwe8kNrWsh/sheFDooM3xDU5SHd4awob
HTFShNJXvBjan0qXhC2lWNzPisjhuvkxwkk3vFmpgIjrtkkbr/PyJhmAYG5zbwYrjmBtEA2p5B23
a1b++XkilcJN0f2r9lSg9As06laxuprxnn5ZR3FLnPyS2wfnNKNWV6ogpbjbVp1Pej2t5fLC68XU
Qwf1u2Z/i+H3h04xrjdGZKziU3DPSJvYNWwDglM6iOiDwLOwc90y2KyRmzzMwzccigNKyi1gA0A3
m8rNFq/aurELRNIlkuKLBkZ1sJpDwGpjSWIjFNtWVIXGRSuBKmMdueA7ER4U8CaAgQMxShc7wY2F
5Z75ptwQdpu4up0VJwBoxSJXTiiNDyjZJJ8kKDjnxMxKYpHz6NLYYHriUsy5mKReilk/HppYTDlb
4AQVS2fRkYSlquTpNFE/17huWNUX5HAYRfmR30by9coO5WvE4ahGGwQfhRkaGyvU4bF96P7RQVHu
Iu6qnG/VyYspXVOE6ic+co2fpS6RHS+26ln3+hRFT1qHH6l3OU7SrwYnoNvrttvKdVE15y7hLN4L
nRPOXPFPUbyElk4xNsHlLgyovKe9Fv7cVX/qp14fPyPQF6SeYRUb1HjZk4KgPnoGudxTNvcNyPYz
Zkgc3E7OoXsxkyvdQnan6bx/7d33Q+T/huGpvrT7of+pMlmFVBx9AwzX9W/+XFeON1ip4hHFx8UJ
HXjeIPbTUWpZgh3Yoe0vv1AK1BQLqxm6TuhyeRHX+7qMTymonn98r+QaLJObjBnnj4mm1JW2i8ZW
3rF12N20ki7rUjiA8jI55LsdkZPmgzGdajgwPaHrNtlOdlwvt6Zu1SYq19wk6OhtQbwmkW0Ng9CX
yibj2NLY7bUHpb2MYt92SozJNJsdVIDNkeNqrftcXTscFMOwuigBP8HQ4PuQGU1cgMF9/lq4oqdn
qeTGl3WlK3D0A0iiWi73t9neISOw6Ie4r+1mrH/LbtgiO7+WIomhY9pGfGpODxRvbPrP3xIJHtA0
AnSk96gJWTYZNtBj4qK35ChSqJNPCwZiT6tOYTo97Q32PKZzff5ehHS/AWe8j7cOokVDwj+jwCRT
PIgeg8FIu3fiXuH6RNyniUFshyBpUktee8hy/d/5LKZPPMj0xW0BVXuTC1a3awpA5n1Ee5VNGEEF
klO4myVawEGaHUAkYq2e0NFY2IGvyVDP6+ucW4VlrD3FKh3bolFsYbhRQx0l9dyvKfj+TeLJLx5x
TpynAWoUz0uzYt7v/NfFVvBX2AsNV8SLzmewCSrZhooARZYdR5HqsP8i3GGbI8WEk8LtijLCp+b0
BiZ4i0w8xSIa4yIYxF9+KJ2DCNDETSi6gi62lyMLPdZIRwQcRpzlqN+jRsp48dBg6RGH9D3y0vyv
fLkZgv8tD6PN3Pdi9mu3ki0kH5DDgmHp9zf5rj+Z2CNKm2nX8wzBs40TyHEa+95lv/6CekuwiIr7
2hh3Q7icojlv/JMfrq5FbYdo9mvdlfBSuXnbQUU6zqdja3Hdp45qgDpHVUEpD5szOKeNZsgRywL6
wLJ2GS6+sgcnbXxFpsY7YgaQQegeCSdOe/H2a1H8bjOWeiM8dt1G2zLCNVoxVkwsB4WIgWh+2WZK
l8i+tb3S9JXSZMOpMNhKuGSrCPAu21wM8BvaDNmOxxIFBo4ye2535tslAXQGQnsMib+QztCRDJQp
HmaRQUhc1rN/DbrojFLPQD5c2Vw4TExevB2wB/YqWhZNKpzkK4R9IYaov/C60TetCkT7tTTcdwWQ
8a/2apRQtfnRPfLmtVvz98jClJgLVu9pLc82Ir2/te6QEszKhAIihmix9hNpRlkvL/psnNu8wjOz
KiHY/1DG1F/+6r7EsxHJ76AMJ27483SGr5QswNhBSnMvto68mj0KdmkIljxP/ZQtD4yF8D5vdiS8
cUwJ3WoIN8KGBxf1HGSJaWHVuS7tVe35o5m/uXvnN8LUi3mba0ArUrJNjrLFMrv2Kd7BuGFZtKxb
PCcGrulU1nQz8UTY9fIFBIKP3AmW2vPVKShrRsmGNiBs4ExVgjSyLuOqOAN39d4cKgPwOO91z1B+
VGikrvLKoN7MXLQVJS+awH4W9RKq1CQD/Xu5xSdqyPmqTpiYhhfixJkJJLhTIirVtbbm+6Oln6E8
Hg7vtu64M2u5nZXxqJYpNmkfVMQoTilFuCEZ7YRVcNYZB+7ossrXWZdXVvmwWF96ZUmmeOh7etfo
TYgi1tq6mFR01ataoidYxJedMYUCmA2OuJQ+sZv48UiDG0FKAIvzGztOzHFePXVJ+qt92c0gG1zF
FunxmLrT7hFSmI4n/tIwSeWQz9+k3IREjBNV/NcudWtQtUJZf1qx3lS5cES/oiv7bz3WaxiPAZL9
aHeyty8IlLugllq4qtavjZL+e5zQt8lPrLi+AUVXBUvHYVk4Dbpbv362hveI8mZrMUVLpbK3m0fN
z+HdNQD/HlEiKrJX9k3YIfUqT7V+c/SWBkRB1vc0MdY/ES9zDuvCjWUPoD04oyUTVLBgnmM/24+u
eeVw7ImUloG2O71i7IuwVWe6Hj1iaym4KM6uY9FYqJc9qEJDG6ZXc687DK2ctomzXRAnC0uHZyWB
hEzZVxtRjT77wQbK1WC1N1D0ciIdHFA6zFlQwmbXAeApx3LIJI6uuF39W5SLxx/L4vPfma+9UfmP
89M37aaba7QAJ5HWpzc3dPBXZFwwrQBV3szZTFpO0gBHZ7J32tfAueRcmVkRPYEwkMyPSaoHmcvI
3bRficFih2LDRePB/1SV0jYOtBdsOKzYKe557fjSoj2FYEgqzONTPpUY1Zrxgb4kojnFEIsI9t1m
dJqvNlKeRhmJ1oqeyeEerpOVT1RfuMgns/cToJ5hzM7zSIXKFmxhBCPfuqGTMHyIV6YWCrKa7Dt/
NE8cWLjOj81bGz1w9SRI41fWnBbK1JIgkQbLeEkgVSIv3QHkNvTAjcOfebCsG+iSYfj16uosXf2M
iWx6gDWDdh66+mJ87SGUeu80+yPQ27wcKIutXddUS0tly8ZZj2vT1vlAJZiNIuwROB6chWGnXuzu
9lZuVFf+EWnOqeoH2UQ10hY9QgwY1nbiZMydPq9XjIvnDGzM/eQXW6CO9jKA+RYIeC3AhJ9T/aoi
fZl2qGvrBjQY2qIO4479DHp3KjS5syNryEEzK4OAjo9h9c2wONUDbsT8t3GsyDHurb/0fAw/gjyG
9Cf2OvSXQxSU2aG7vnxwV8wQ8SrmfIK64GDplIheNICO5EaaxgvVOew71FNljp+xqyqzdFbyoa4/
pkZIHhyQ5wd5eelLIKS5eNnLVMwbU1HqiwDWR2wmbT4Fxi336HC5Bev5b7hbpyYzE7ZSGCbgRHcB
LOmDPjZEXCvTc7KtyLekYB141yGZsIpsY2fjGDswW3/GHW8OcwmQ6EKqT3m3Hemp+tK+W45SkwGs
a2xSJLAqtrcB0UwtMOYThOKX+rIpoDqUgRSlY2WM/S3ZUd3JVl6vIsdchgaZ74XXipcP5byCNRXO
J0uj6buIsntWQbuYN4MYackU4fJTV9Nz6RwzkqA+5L5gzakXY8KxFP+mCzFm9LbyfR+Z21/GwCGy
xvDjlAES8yicWnGR+Wrh61E9Qm7gIeiyeoC2980naQ/PXRSsMZFkLE2uqNivZbruphxCSQEnQt41
Fz56dnhA9OnViC1pQ+5pok8uj0uGNhx+4mNnw6fac6RvO8/gt+3QWVTN9tNLntpFzQBzn8vkULMK
3G8K7YBrQH4A0lWEDpKNeTzvKa6rCmPrBm9t/LnZwrXRwoDmzhXpy84reMOUDztFGFQGsaHOrB7a
2o2pdresN47qfjOthIRG7WJnmWr/GyFO1rJG9QPZC3cHnX3CCyma4m7XTRdz612GfYrRgAXyp6f9
1Xgj+SWdXd3499vSOmAcmifGsnKjfeKQBJNC9X8Cv2VvoY/+JocT9ipFFXoP1SSjfaeQj4RTGY3z
jKaq7J7Rix2WhMeqhs72UW6JR45ofeFuY7ligoDvxA2TMAc2i7DpFxBJALhC6SsZWpHuV1udk98F
sjhE23NskwU0j3fBQ/7YPowttyD+be74SQkcXeeROWjNYQ3/5poqVPA8f5ZezMy4temcuw9IIL9S
lU3Zh+h36sm/K9WocE7lUHjn9o4aiImOOaEjeIUQPS/nZonbLYqEdEWHdLxC1cGHy0a17CP1v1kJ
7RP6an+ujtpzck0kavuBPO4sslQj5kRNiw052V821yqDYh7t/hB5qquHrJjNj1FVPI1iTD9xnCGi
GlxgQUyXiNGTw2OQfa4jxtcCLSCaLDBiW8GxMmPiaaypGBYfv/kpm9yRxKRJL2/09zmOH6Epd/Qt
cUqfJXKkJszScaOiOm4L3f7SEzjT4OgC0zipHh9/ryPNUI07YjF+lxhCK0OGUjUnuUAgt3JMZ1p4
EenCqTasiRLMFEvGHa66iShPNKmp7dC92xoD1XqvuZ1aQdjbjAlfkKinUzV4C0Qq1D3F9nyUwnyS
SUTkqBaBhBMa6bvDmnl+zH147sna2aR6/9gTUagtZTVyKndB0ZuKcx0GWMnj2fvtSLOzy/rbDx9g
FvRrO4GEt1e+EE+MM5oFB7YgEur1VS7x70zLHaN/6a8mAJJX95Qq0/PPq3n5MWvLmjAvXTjKepOm
wAoPUjtEOyEwZVMtl0H0kY2OTPo2YgSNKS9EUNoWGPlznqaWAU7xXX9ihiwEHdNyof7GXy9gHr9v
Eljm60bjsS1SqxBUdVGa8aKyDltcO7Y7xNEFks9OHtkniB25kCLUkLbZC2KBlAj/0+77zDHaHxPW
YaPEL5NKv6Ro47hvEFgi8H3qc04GmmB5b+YqjKHThI5fvrQHXThWsKP0wlMsbkneE/1rzkqQCiQw
6OqBptdhuv9yl9zj3TRCTmCD0b2Y/zyYFuk1zjjKX1kMx71sKJfGnWDAdZTp1EIBVxkdy2jZgnnA
264fKUYmvsUGDukKkuxiXptrlo82j6lPOosi03LDveZ3gTx4yLPi6wvuuON3NIv+ULOf3UC78Qwk
ORxcj/Y5kdYjGfvFExC7NUDg0ax6b3105jrQ5l5ny4a1y+YiiHKCcww7gyYmASyN6SpnuZJuKEqx
c83UyLzL6bWjuoCHaYRh7gn/PF/9OAROjiNEDTLCfiywqjp4kxrM4wKjiSDP4RrdIq3X1DsH9T7m
1vE1jq01iXlACYqnH+z9F7nM66ZKf8FCExSOJ4TyzZXZpoRAvsUXL6RYXAo6PpAmSvCORfwujkRQ
AR+tCic3YsbtUUE7d+70AvV0OenN8wPYfRsikCwkcWeTx7mn/T+za9pMm3QdjpIVCNyjKI/FdpkP
1sRLqmWCp1Nxuf7FpiHZlCUlEpNQCtHuFP5gp3w3iEEdpSvedvUYHhxXMlNp9DxfwZ3japRJFjkc
v1KB/vBMJascso1FoaxPI1TTHoe/aCfVf8GwHX62i63Q1azkm2r2ckKel1PExxl4rN84uVfBWuFx
YA+RXBNptE9RlN/oYcQ9fobzi19TuJtYGHOGm6g2t6rzvDGaljyP7WzkLewu8iZfpuqgDm6ekL78
H+wYRNAuO+I9Xd8R9sIA0zmFxw5ogn7PsvinD7nSRabUyL7CyRfxIoPP9OK0FXDFc686YUc8H6+X
LqxFaaX3c6Eralhtw0aExZcMF4oKWx+pgerZH/y+UqyC56hwThewLymrmiYelzAbi8253heCNDKn
/QPToVMI5hYSNWhX2JyWDbpMADleVzbWnbeP1SS8VD1CH4dicEjzjm/m3z1hSnl7i8/e8I5ckTjb
/qAg1f/fCshWF39GG74cRuT2vd6oO0DGtEgkkclL2uZYRHDjL2CZuU7B1IwmcPoc+AeoUGjN8agc
NmNJt49eMeoMV2aaM01fHXeaGtO/ko+Uc3FoAe5oOa9IP+Dz6rG03EdV9iOOlUliTPqRrr1KTEIz
Mt6zIiXUU/Sfi3CMAZyARf0usfHw77Rkteg+ag3kzY7ixOjLjDVoDDhlxyQRNG/ngWUikvEM/GZN
RHR0DDAjxkm1k0iUdmcHI9CS5bpm18AemaPzDYb9atNRREk0xh/bHQATBo+NAqa3uiOeE6slGry5
nTHwys3mU20CLG7nIFEvGM7SCkDoLZ76nFukQz3JrnKVpYkHZI3wUlP5te/+GBBHYVvMkVXSiRia
+8Af9YYhFBkEPBj8UcU+uL1dkpkRL5AEpLCCMm/NKLnUZjuJ8gjlJNlOsLiHJHqYescbTJtCZL+O
c3clRT0L/2z6SuyBiQ9yMD3rlfQ7EzJKT1ToeZA/GGm4N691vDiX80/yXPgoPeda5I50ZWT6853W
8HX5htuWEEfaRhxNJWkcuujqG5c6xS7GDEW7u8b6cXfjfxoXvRGyiKL6T7+w6QiT1VDAeoLS7T1Z
zFmCXdhA1ywwvtLGx9RX2I1dGkEQrnjx8zylI6fAdmCmL5uRF6rs5fsiVoZdtHleqVq/KeWSosZ5
ggK4uvAAujZCT4LP2kgkUY66neFDyP8hVa2uDWd2AckFrZ9rPK+jJj1HOpLDq4YOFhk9okn72204
qeefc3Q/4R3lLOJnBTxZ+nDVHa6fxnXH+cbMlmLuU15yP2OFyUYD9tIzAnSfTSLsb4b+4jF6Ehu9
JI2VoGW4mZs8SFXU1D/ytGcVWupAOrUPPYYG8YCuz2CMCbvzRZxjcnW3CHZyo8EUOQmYG02GYhpX
Pm9w16mipXITA0mpPMstSViJd0oSNUyAhodGfHt74F3AEtuIkQB6DLQpZYPqk4Gcq5pf/u2hV6XO
BBr2M7mxTB4MxofChOqF8UzORQWTHRVYppqD4dJZW/ZWbYgfFz0QnFu/r7RMOaSFOVUbol8AqZ2M
ta3Ux+nvUnFSdZSmNppkOmsEsYr2EL+dJb4OCvXKsvA5Qj0rK/k5XWxvB+H8Uoq/yPE0YctnVtdo
nYg3IMshYUYkQkj1S89UXN21eP+zQU84BAG320VGCkBOkKDeRRO2pmOntxW7vXVURpyBYLcogdUT
LvEzjN+4vlqUkeI+lssWu5+Ym6GT6+PbjUsGIMZD2dLtjDqoQkRtXGgNXKKEXWiobZCUK/p7oQ6h
K1Ot0dx46EAGhwW00+d/GBD6rTGpRt4Yb9xXkp8B89UEMghjLioevOiqB29eEtbytqR08+hF71Cg
rYyLBQ9n2Pmz5TorkrUGT42ATfefKtQQ+MZn1zKQ8IiFuplRK39n+IJZWNP8NA9iNaUmtXHwCFVN
Z4wqJEMAJhCIdSDNFd2laSUY4Pahl6U6NcVqebGTdfDNy9WvjVFKeg2QROpT+pyiE/vtWtygxw22
mtvd/reDUAY4zTIqmfnj4bSVLGrxDoAU0auh7qzamnWcNWQ76xEwOz6wlr1BWc5ZgxvxyhXBWmsc
HJlyvWYAKiJpchbxtuRS3Plr4kdecU9AOh4MT6OUSv/2mU0YuYTXjLjrjUnE/awI+p/VY5tJDI1H
z08QK6HjkMjF/TS2ucAPqV0if5AHZKSlaRUXWqH45KrRGoS8Zhpurk4i4+qGv8iEfKm5aV9Xd0y4
OMsfOibeEUNxc5kQdN6WKb0CH14Q2vUcApUzi0L3KCfNyPK3WFaofaFPcE44tT1xDinf5o6bmDMF
xXabWvoHf+CRwiwKgtQXEW1tjKQCXHDK02yMsipXV6qcwAaX4YXDDs3IhmwoY5s9NDRIBk9LU3UO
V3s0UXdy+qhm0/Q9Gekq1IYJLiLFG6hETMjfjakheCifVQB92+4GGYprOijtVP5tVl7bQ1mJC47n
Y8EhaVBkaFeHJqrVWbhoQRoDwTB5PjDmK2h9Drt8ZkkiNNXkfABpUXIAacF+zcPZ6oKVi14i+r2e
iXk4OSIkBlzgzWb57SJ3kCTDGyOR5mbrKHEdqAv0xqfuZN12dbVS6mAAsEnyAkNA737m7/hwKBuM
Ss2XI1YmZstV9QtqPsC7PrOYRGNCAZX72lddhdmZXuW3/PItlF//Nn67RwpoJJ8yEIeBlplQ+PYd
m+V8M+ZtZFNL5asSRJ+upAh56rUjsoX+rtX6I7u2jU+hR5WOIRWDIt46QmQ6g4jZn7/YnVqmH14v
UyqBLZM/077UCs4NttVXqVMbHrS7ANDQ1V7DGDMLFJt8WryQXKBP9yNvHx2vG6ihHUZdFoatSQ0H
KyclZemUz2jERWWuo5h9TG9vh1LVPP8QFyYdPYO44ics0y3dzFJVKT97GR434Lo8e8bqV7vBtUPO
ULsaxBvOfowpGpdzxnKPI8yLIABL0i61IqM9JxZtX7uDVUjnKiZbifDABuqFCcL0hVkSDLpjErnW
/Tu4j71unPflkIAzD6K6ODPxOekVlbR8mKAS+YKKe6aYW4dBbOzo7WJdxpmpR2QwEPHvBcT7vv/c
cqfDZQNgr70ZW478tl+UcsSqG1odH/f2eRmf+T1x5lAVeLKyE7e8raBpa8SrQP7g4smZ8UCCY8xN
LDeS0/Nmm2xF/QNgpeCXvzK3vY6+P4pfeTMovbNK+kJQEr44Yie5SA0EaOHmsm+MAA+zYkWN6yI3
cGXrA9A0ZL2NL/+tvdYfq2XU2Eo8r2s7qEr0p27jcITzRYJaja0aYzVt9DBmi6l1/kzDk9I04Kns
WDSHdxNtvXCnoDVczWdMu14tZhD7WtRencdPsZAiub0KpIGbkwO4ofwfXbAjjRF5j1O8qZ6uMBjJ
eLPGKyljqtrM7/ttiwWTpk3b2MDQDVnLtFoIQL/c4lzFKGJrbU2Q8mCl2RGMKUu/qB6SYwayGtbX
Nw7XPyImsMmrNcfpAc6ibGlvXAXshNylfrpPxUMJ4Seh+fRz9djx8DYsKJPRRagz4jwYof9rCOFa
3e50eiI1kzK2ivGZqufJxYk0+6oXrrMKVfDmvllGmqjuuXtGndFFfuOeMZunj8i1+aEcJGt6gnM6
NqXz9pNzcTaSc/WrKPgGBd4K5dgCRMUuGJuDRTBxn8uK/M85fHke+K+PMArNkQIJnaZiDZYff1oU
eSpcqVNmPhaoC1APEnOZck8tthews526A1ZGAeD1cQ7HKfrqzxpzuYj4sgqyHHMaFI0vYdbzsbws
jncf+xJglmgsfDUUtLXNj9ej87U5eRNI8jNG6zwE8kB7p6jAVwFkQuNbrlzh/vjs3HrhGB16nm2H
j2/yyPLHSDU+1nCYa47N2xroTrpsYpV/nZwa1PF5WBj+gsoRYmiItD2+yRKXzunYGYKL3YbI88eu
GziECiLEOYG1bK8qc6h0TlwF7Uka+28oSU1249BPc4SX5Mccnx3ndJ7dqoDUQMV2MCbAP7kVBAOD
G13xqUUa8bCJIeBmUtnE4791e1x+6oS7MFlmk0fbJKsPxQJFM82GGbVo2zyQjh2nNqlXcBWzDmK9
YXAJ1VPGwvCsvOrxFx0KLBrdEIhEccPpWa6sq9xAsFJMcVJB/7FlOtyFQC23ULER3PFjAmH+tYo4
P3pTE7f5RmwFIm+fZq9cmEZ78pbdWQTQlAShnU4rpnheZ6FMdiVBwj1Y/DSPUBDep62T7wFrwZbX
kY1qBQhF5XWtr8a/vIxae4Cgt1q8AsAHeV6IgA29DMF2OlAtXNAgchvTXWyutrb3BnDvCW4fpiPa
8440GLS1gRMpNlQv35Q9rjT1tx0yVhgHhha2/sSZp8YrTiObAhRfv9frhdRV/fL0E2iTvrj+BlnX
YhG+88ShDJA1iWPArZJB0b2Wqle2kdiJXhUpp1tsAa0JzKkw5krqNlssgDdWBOXSVTIoU1THCveI
C2K4vcOqcQil9RbSwKhbbKlTT+Fu15f1J9ni5d35wrvD/Tn9U1Z+1FuQ061jJcQA7DdYB1nbzGyy
NdDdgwgt75kKEZJkiYCggswZFQpcTuvqx5ETdzbEMWTWeonfFJ+EBPz4t39m40ajQAUzi8kogi2F
4lajmQTp4eT86zloO8NkmqMYxZdN4UbcC2tMm+FmoBcfbgfPV8SZodUMh+TyRX9CaBLPYP5CrEjL
j/MicXvaQQDcYu/A25Ni06LlAUMomqyHnvTyohQrap8YGJPm6RB52BEBoiWFQ16UuawJxUts7TjX
1yjW65V4Y563FXKcxG7knBeuwwER1M7/f1CoTen2STcZqbYyq6mdu5K3sSdq2avhgZu4MxYffVqI
rwCNAJJlFGjm4DiX0mSTuumysMF+8QTyXtmN4AWHlQ9xAuZ36QiyJqMF+1iUunbPR7rfFcZ4Wezy
8pae/HlkTZn20qfh8OXDkWr58g06A3sGyN98iYSZUOBs2iP/XXfhCtt07U3Ra+pmN1aTMhsPAyau
5rNC0BnCly9p4YnCgWN7HKJMV/uCoodDFit4gGNCc8ZNeFJkB7A6F4u2iy0nQSFV+nKYmfUO3+PW
VCH9ai7AXs2sxxKPUvJOxDSiz1DYcIXLGB5wtY/4/1hONzSEStQ4kkALTh074pIMDydOZpYCRfw/
gvQuYhSz+XEXbFWHgcZrP4PC9mnd8XBpSejMv7I601CniAAv3kXQEWxFTDH4gul58LEA/3zKlzti
608B8HXmWNMFp6+Oni/gKTpUtaI+5PY8MavNa8HJ3b23Y38Zuq7VYu5TixbBajsPBcfqX1gOaZcT
Jqg8cCsVRBhWIphWa4aGUHfuvSgM3o+Lrouh+3/hNFtYDuMHeSLrNGJGz8FkW7Nl5yRA2P4z0A1U
7/uRb+/BHjY8SXEZtXhgCC3aPDHSnxtSBoqVQhPmfIzZZVjL3cBWbhMxeTV/qmGcSlCsnvU9XZcB
dj98mUX1uIp7KsIWgoxQBCCTNplyYMEXCqBGVEexKGNtp6ddlu4oxqO+S8A9wJPsO3EI22PBaSXW
9LRUc6LneH9areBAz6rQb6Mxlnp0ggpX4TgtBtMQwjDMateAmg4m/PEs/EDYlSVwuJ60VwPGH0vi
P1CwozWR7vzAmon1o0x5v8D8au1RmpzJppAxBTn3cy2F8Iw+i00wrIOo67A+lFLcV7SY9rxmYAS8
dnQpT5LLwJfTboMuDTLMo0UlKDhSJBO79qX8gLLCWvk9i04QfjoNtpy2Eb5ftVCBZFjXufoCN4PB
ZfH4IPzclNQ26XjbG3e1KSh/4t07zMc1BpJTPk2rfhdNwXFiJ66XRyHxlYxxitQRlXfZBwVZOWEm
ZMX9RI+L56hIHVxe6fFuRljHKZOl7aVzU405J1murypjiccsq2xVq8TAnch4sepgqK2P2UYm6XB6
MG4xs4IQWJi8T346u/3MiDNHGFCH6fedb2Ozb2ASYeQ9Zebn4nARPdwMG7y1ptcLCnieeRGsR1iH
aGwyS7AwaG1+irUQYJXQkcpmDgzsPpQB4VjOam7CNGiLFx92JjT0qdWArbG07cGxkzR6zhAMq1uH
CPNvKPIgA8hGRGk/YpMmAjVWmLwCiePGKGPoi7JKyv3OWYy5dKrZCQ0KyeSTmAGyG19n2XZBxYH9
U8oPeFwIjpeFbGY0k6/H64XvpIUY5hawzHWLCrli/ql2ImSQOR7hUWx8QjV2JN93zwrZTQCvm6ux
L8Cr3Ya53EraXIAMdXcifKlahh95iaSuYH/4AwJpWuyqTkL4yibdacmeKt69ImhH7D3W2M0Yp4t4
TAseGXlP6Fo5Qm/hiHIuxT24zGTKaUeZyIctEyzoDfuwWWCXU98MJ1XjkI9ry6tJGBa7zn5INHwV
KheVlUVD+Q6dvf7/h9UIPkW5zwY7ZySNxf2/Y5Cj0IOjCXK8PHxYxN7D5Fl1P808+YB3HYl4sayD
Ib8E5nPybc40ZjF1LL8iJV1e6ghJtpeIIGPUeDwvZXt5+OOl/r2Qr9PsT03rzdOfmegGjKOPsy53
+qmnkOUoNoGYhdKesezzQd8afY5T3gAUefsvicsfoJUlpJx7XvyOrcP6jmNgy8kFrzZTWZ11kPLy
iY+OKqnVVExz56nY67uaS45j0jeckvE6gDx1rNsxBjuKFe9edXimEYOKndonWj7i9NtsGyaqLfwL
RcHBgpEjn8O7LmH0DZAW1RU2v8BQx9Jcwckkg9F3mrMuoNGAUod48KUPQ6NJBmKCKGBWtrcCZvXq
5VPSw6gDVBHbGXuKljkW93jX5z0l7BKX/wy/jYu5V2ws51uofXPDxg0KEWPfOvG4WJpL1n241OPF
4MZNxxaUNI2PnX/X0/NNI6+k1fOzIy0BfEndVBqxLSd/3NND9Jy3rI5rDZX87SJ0lfpHv3/FTwpm
aCjsVa3nRz9umghom1q2D7meldWNLd8S3AIXYwb81Joo/jyDu1iiM7gRK5nVCQDVB9CNwb+XwDdA
Mj6WhNAYph6LGjcxFHxdnKvGyzeklTchyInrCRoHUBymDPdPg4teP99zuhDwl1dhQzbo33cXCMt+
yL8X9D8VxjUXtsOnEy/oEo6sNg/j7C4U5SFZlho3cfjSzUv/lTzu8Ud5I5oRYX5nhO2i0XlW662O
zoGlEiWJI5Fcut/Jo0atbS5M9IQyp4Vi+EWmjslSnYMJ/VFaD5ROCx5mGj5/8/1ZnPXiY+HmUOgv
DQgEqdkKGEhQJKxRl5OddYZBZQ2nY6Yc2vCNhaPtRELHytgM37EDdT+0CWRRjHp2MRrkaTkc6H+N
8XFOLxmwWr+slmlouoQJxKtPZ4Vr3IuNoI2ApSY9E5WwPl0WPOQa8nIHKnHsZGxwOKXW0VubopdI
TCaIMK4uc+m6/LPhOlRW7FO9PvVuJHmCBLrVJQWvrYu+ePpICBfoXrM5PsUch6UG1PpaBhADTqRy
ip6hEO5Gm6JVx0h2So2vnCjMSXfchOPUQWUH9xydDr8DoY/RwUW9kuQT7x+bkuWaajuBBE9WtkCz
cfBUJRSbvIVlI5jV7+JpduOia7LgzzBdAkaQdDhD7MtSr+DvbOPSfKtYmTsLzkZ8upVDZiPD0woo
iY0I8o1gI/UYI80DDmIg6dqovBJHYTxJAyILaC7xugR8bQlmQhw38f7v6Vy1Kzfa3S/NBc8IRe5c
xZvUttqTUwXnSrcWN5iAuzUHd5DQjcqbyIVeCDA3pUMLOfkZPqd8DTHttl6H8YD6tFAfZU9oTwV3
/VGF0FK+gIp09jscBziplG+oMXSULcFTnBl6QPQ9vLeVYl0USLjvxqGVrDiDPykFQ0RuEyVDjmfN
BR0swLjk+hBWJ12CIzAKmyK5/+J/4UL3/fBGqZ8nyjnnAxtZdL2ttf2Jij2vqyyjl0pjDVTPnJ36
yGY1pe4FQY20kARYosEbvo2pbEmzNBhk+cOgvLAmg2jWHZBwDw455Xqb2IM5InhIiHvn2peAMsye
eG+of+DLg+2wBeDL6R8KIjpettPOsPD/xI5SezGx0469dyp7LpqkYwSG529Jhr12GQJct7b8R31V
KSqd8WWoZyZaW/3Tua4kL6p9GDPkrFMOpmC31MFBh6qDhlJNl/EfZkJEWCvXEiYljPb9oY48Jx86
Hm8gUiSCIC7T+xb62l67zpeNR1ENMh1l6IfJ7NbFaETvoUgPDg76l2KDJxS/2eFC2g2m5+tAdA6o
w2LhcZuntmU81TlWLSQuTQ8eJ7MBLlhOUyv8KezO+NBV1ld/24yaqsGGfu+npenc12MMaY8yvIQO
1ijZhKph4JfkLCtxypBtXZ0xbML5vZxDtxAYcfsGSnye7X1bMg9OQumWIfw4n2D+9YYgXUT6cTlF
VZPAJyhdaE/56gOOfzoiU5W/lG4fTERXadtuUsTEK2wouxScyKSRjfB2k979DCD2tJl8ecQcKger
ZKwb/42Z6ekQZWG8ePR+HS3i1hoYiV//AXWK6vfFT4K3OC9L6ggzH9WNMvbaX6FztRT/16KUsbkv
/7vZyFMcWbVAJT3EfNPEhnI27jJnBvDfhRaKQSoUO6ROyhdJsPA6qHeCLN4He01I3TDqMERIslje
G9avrz6oHUsaeKUy9dV7+sMKlRcJ4/SayY0ckjAQq9OjVi0HbsT7czxeGhW6unyhM3sTnIk7G27G
Jc1ackq9dBMpkcjnA4HKWeNjr05hpR77gMPbZ9gvfR0AGwtPKtmy2H6Bpqs/iRd1EZsxSv9FzD+P
2VsZ9aSYAoqNHSa+/y2adOjYxp2gSdfcjb16poI+l/HaHkXkO5BMRSX7TyHZQMQ/90JJOdO/aGsw
eZftP1qVSmRqfhvyA/lEaRYRUcRh+3VClUw5C0DpkeR/wrwjkmOfDijgRfBJxC83BVSra1OpgjD0
hv+NHbkv6ONd1ducSAXDlV42416lGvgBr79OB91DvYaVBnTX10H62a068jSXL21Ujf7JmLvxYz2p
DHWPOzWg55O/OC+TvgkmKjUvsc6BXgElNTMc9Xzw5cZ3LN2NCC5EBAIi+pLN8TXXZd5ps+YFLtLd
ZoCn4+u5CKZktuGwfLjxoj6Yizod1emNxcrCU7Q6t1UWfaiLMvH/dGx6jJGE6t6GM6zoEv6UXJEd
eVnaJZT7LneWizPcQEEmOBjd9eAk8mjYURzCFQoMuOTI1asFWjhdmI561BR6AAXlWVa+jFKakJwt
A9yW/e6OlpsHjIaPONaJC3VKpIg9Lxb82jwFa+EnZtVtDQgh19lCKUspLOgAtFqBwLwRvFS7filE
9liOYggL3xp/LHUVIK//JN1N2CU0/zRRiZGY/kP2Qv9uqG3afdydlZsJ6+aglK+oN/r0WWL9wPeS
HAAoU2KO7UTjZwJ+j3knNOssxuq3C67AkkmWYzvIBA0Pk6qF9hTYNBTycnDceCahcQjPjdnWVx82
GFtmMcoKY9DobOK90csAzeOivzC6F6yehxP2De9PkEH1sWGXFxWW0H7DRehRhTpgD+/4QBzpAoxu
FLVRWVO1ZVGr6/kSEJ9BvEMUI4zquEOiSNHfTWw2w31P94tVij6+xHpsZl/JiWMtkdFCF9t8DdFK
3e7d1dm6X/tH9t4I0PzKhdjA/kfIy0/nIKGu/yf1P3bLul+UYDHJyjD8icT7mNJrDQO0oWLShNTy
5Zu/I7XVDu110Lw91t/QyTv5z7ref6tIfxWuMM7+2ddCE5Q1viQp2af5DEV4WL0CIOH+ZhqAeN+D
vDh3pEkHv6U3931HEw8KKaMKa113rVfIYQ4hF5gvtyfRmnNBnq7J91ugR7KvsFcpTga9eytSXEsB
9Wx4Wx92JkZP9I5TTl/wLppaK+wutXpij4NDqhEFNosbqA4FEPI6m97G7L2vNX6WkfPJG8reJnkW
UhMPHPlmkpXOkHBTd/5ef0DssKa+Fe0uRvD+F7wjwU3E4JjVRL2K1NPZn7p1pReH+X/ZrFHV68PS
cxaTmyfqQoQdYYSQW+1jf/dS2I5emkDjNU/bseTZXIjEtK4FrLUeLCwbsQ6nD6jdfU7arkyff2uv
eJZnXm5o9F9nRPXwe3Ezas+bz59YcoJB7Wr6AAKXhJwA83S0LecGQ70jqL6nXOjdQuM3EADQqUzT
wwtiGo+fNV7pyHQILq1/8IuvS/YYfI41fhEG3TluSu51tL/Cyn5SHnIlqGYyqapWzt3/oZdkFrDE
FiIGOhKTi7CTWZaQlvUEnU0WXDV+JWinMC4CqjGv9KnDRwrsIP7iySvw4D2W+zLrRo+r9wn9eWtE
8rPD/PQp8ZA4b4Xlx/0KOZ/G6BbfoaZ5xczCC1nkzji7hPgTNnt/PzqVjwwzaliYvMcIjCEDb5Ap
iULgqA/ONKLGbSDGIOAnX14n5GHrv9mx63tVggdadsBIRqOPV5T+Fa7p059V+TU3ReXHkRiZqaLh
JI+UN7zkWN6xoTCViXaYtAepZI4vlRzCHQuARXEcDaqU4fHRFBl58KTnvbp2cO/K3WHEyq65bgwh
6fa3THslQ0Q6IyGmFUtK1qV/zP6emDym/AVbZNq8cJx2xE+/cUhKiyyCTZxwra3/EmjL6H6/JjNJ
UX8JrMsS7dv0PYyryeZkNdfRh21gpJgzQQszIPUB0UpHhVB+JrMNdNaA3/bxO+cyvJENLhQ5h9vR
6Ke9qdWsOOnMizt0K5BY5Odi0syvoaKIEeNkTo2/2/HL8JpLJKF5r787lW6LjtvL1doKDfFj/fZN
mmCmxiStTR44BXczmpfdb+rqd1/IQapxZZSqb9N2XojFLqn8KDcJca/Zd6OM4HPGz2VC0ckqoGOX
eg+9cpqN83cKwBkfbwzeTm6SinoLQkHCPlgSkaygBegdoM8qqQ7kkVb6NC+6pWdUgXW9hiDGlF3p
qn3eVSJ+6ETu6qSIG9wSRwc15FrpLWBXnOsNVhWKiOtzFKgr8iDiWhMwYy4YeowsB0iPwrQDAw5Q
tvXKM63XzgbjKdIIWZgr/99Yk/1ey4BbSt2d4puPRM0UcWzVJrAflXNCJxW2TJuPq5CV1hlTWZR5
L7WefHbZjyCIt700u4QX9jtnCCJq4Ys+vkLu1et1FLaQOZHhLPpZDGrZMz4tO0m1PSuLsPSTpzr4
scjJCOM8pFIbBnEnKxV0Cg5WrA4IduHxtE50O3475/s5O7pTum9cAf0No+I5GhB6ls6kARMobwC7
vafwpsUkjptzBlzHLV3BPbFsxD5K0cK/VslQIOEfJktURID4kgwTLubmWOSThupHje7UOxps0L+M
SnzCyq7cFbPoeKCKt/4x9EKmXJuIWG8f6sn5Wnu5PN3VksvlGp3cg9liBW3NjPWWI8LMs7iaGeFP
0hJV2dwNkCGt9v07EUAU/6jvva5XDHh89ii4wV389r17xW6zXDSawZu9b1PzjTb84zvwNtkQG/l8
4Bk0L6GulaTRBsbUToYEJhqiJ/MOePzCygGMy1K8Bv4rZgM/X0TQKIZbsn46JQeXSEHPitfrfnZB
BEMgLd0O+WGRO/JvAbt+mnSW9A76Hu+qQXPa+l3I4Ag9iTj+bHdRBb7rN7HX0K88I0yTrCE6nNVk
AqjdXiun6SoOLU3uB6MzkJBj8jejdWCAGMHs54Npxk4+aUBHkb8J+wUooZwNMm45lY6aYF9PzIJx
vw6PPNd8mB5jJFTefQf79K5Q5ZIuWie1zDOzqRTPqFF16sYx2hB5LigyHeucSsZqakrdO9suzvzS
5lL6eMV/3E1p2a4R/CxkOGL+15sF/+kaqH1Ztgk3xuI0hpEp53MVW0saknwyoEYroi0hUykWe7w7
Jo2eCIZjokYB6lEyBg9TFOA/JjvvLUTigLEfpNXvccabiCsWPJdY8EODhLqFpHHX3wPzs6Ox2yPg
j3qgEqrQjGORlgiJCzmY7XsBFvzZsA1SgN6/iHnNdlj9wCuZsJZPbQRLr5Lhut1HtfVmkCH8fXKA
mNywLels1StKR4hrhZ0fBv0njucU8lMgKrOhmZqvhm3vS46c3HT7yRP9hzFKHhuDuVBptAUt2Hd9
fe9ykmzBczfHVFNv489VxdLApKCs+MhdzfuyF2wfurGjRjYy3Q8qPmCFSmM0K5smvIP9ViOk2NWw
p8tbqCpgNjI90t5hCTvtUIW+Q0xME95wfnEinpw1Dm9AiC1bCrLwto4VCpceb32JdFLCCItCVjBz
xrVFAJ00q4HvXSF0HjSxlN6YBmpEw/FVI+iYqSWaKAh+PzTj/c7yl+AS1QF1g7USggmtUfqTlQPD
VTsaZ3/WgPB+yPZAqOBwkUBSGxz0dTaVlnb0g7L2U9B6YS23x9QawHbln9A8GZd/8Fa8ZGbYOeJS
LxYG0Ke/MXXpqQ+S1rUTTthmDr6qXgCtrBZo2nCVvIQUNggx/RJtqZFzS9yff0oCtdObFRv4rjW5
fXldTIsVGhpSm0XCJaft3+gM1ZMV7NW/zwNF/WOcj8KHzEt3p69ZqLaf0DY3JetsrbTwSV3Yvst0
PKSdYkoEOEVPOorX44MTVeaR10yMgC4HwihNpgH0UJ9lFAz2yQu14MpQdInTe1EdEJFUrN8/FRpR
Hd7y+JOjoPDbmMbFh9anSi+jcpLVoiqYD//JS0QlHaJMbXbjWYOQvai54eLuiW3Cg6jZfjOeGPsW
Mp9QcGXCE6glz5rKfTeBx6S+Ftvk2hF2bxUZOnioVo8cKwFhT+AQFHQXLLLk/8BK1FLsBQmc9Kkk
tJN7ykrN4Cp0TA+zrF1eBpf+Y6dMwKjYPPpIaUh3Ilofs2griHtCMzLnauh/2v57TC1ZDLts7Gg+
VEPlXCquOYihqYNTzL9Ysvygt/U79q+9WzwEiND9PCwJFBqL9Q1Nbl+h5ExnFx7rzfkVIhAjrH12
Bkw+0vwtAWCybQ3vqvI+aVxhuL3mAWLso+zVUucBMttxrGS/g2gv7bOkOd6DzVDkG6nsB2JjmKMP
S6AW+STBJLtyMtV+7G8ueyrbBEwQtalmI9+5OThVGpsgtyqhhMiJ5iLTeNl/V3jZF+HaeVu97AyB
3jk2ZJxSZNa9j01Ac+ckKRh+u5G5w+kRlqvlpUeopkpBBkcAcobQ/5KcNBXihcZShc1nhVErrMYp
e+USihJAj3mJzpDkn0ZV0pGPhc131CPjJ9OERRB/Yf4RSsWSY+15SXzT4GsqwoPNHZ8RisPxq2Xh
U3RJYc89EUc1/KATGTNII0BXdhylXcYEQdm2ZGaNRJvaQBCoTWbYKS3/Wj+owJxWgYJkxrBz5o7u
qCBE18Q+RXURNaZHTVPDlQP6x3+dV3YS0w2GppuuWX4lIQoveCJyzGs7Bx06D5zx0802RO/GIV6Q
dbtmnWqhd0TXusGOyi0dSavaGsPKKPm69vKzNZ507vWy+tIHQhedoUXtHiXu8V9J/vWsIzTcedrP
SvOu7R8e8dMepUhQrtdCeSdARel8QTKQVYKY4ivw9m7ZJqEFKjGot/0eG2NWWSYjeiNj3Y3ENSy1
692DkC7BZojyPP/Z6G7BoLov/5phfLKOAo3LfP0axBNDl1z5a5oQcssYKNQGEZA1f4X0865+h8Bh
bHI1JmQC4uuozVw2/9rwh8gLkWI53cZRjb9tXgBij6AYqoLntxhPGHCO+rZ/KrVRtogOFQgXMFhs
t6qfQWbukZMQZYncLqO2WA0+oNFEXD3CJfoOmbRo7QJ1RokqGFCbXJ2oxTBlOnoQ6st3efGqEV1b
7SdH5mGcpMW0zx9f8+SggIw8wUKK0mHIzc0aLYPpe+n0+pkRiXUFu6vWrbu9QzVO0VEi5Lsep1LT
e1tyxYhuIJz4ChTV6o5H5fPdAbh12ArhCmkySDlytCfhTdvlRv3qFJ66ccykdA7XOiBdBhJv6UG+
omaEcMvSOCOmtbbum8BB3vCv4PArvemLQYC17G7o7uu5AgTeizM4zWbf1hI6B8C2YgF9mYRipWw+
wOgkGXhDDJZb6jOxr6HeEi+Jb3pMv1ujZYQiQq8aAXDleOIe4U6rrt6PVniWtc/UdDzpv+7R4HRO
OwTZQy7MyQmcTTefpxIjJyOLHFl5hl29+eXrQSk7xEZ/vFywDSOm6y5uMRmkTaZeBHqCyHbuUfej
r4DWn172c2LYJc6dIyS6GAzRjF8hI/62zpQ1VXztPvcEkCr3zvALUZx08Svs33lrHDkspQCTtaD4
/Mvj/jk7ucnYe4X36Vf5OVxGz9WlJfDmI2Ih6gQh0sTo/4YF2fL0h7yViu1dQJBqdgv4VHrnvkL6
86llIbhlIvApbJStJomcqlGemzaHmgF7KZWS9aLiBs9x6KgzNwLXG6djebxwV8JiUBfbMl1G01Bk
31s4T7zconYkmOqZmyQWKhBOSHVlgxgmfLfMv1oOq1et3kiuB9lVNngMdYr0riakRMcibNcRJ85x
fd5uoshIH2b9sShz4uUK227RxoCW3Jr16LACj1JrOTN8EuO1J1t1dGxVRKAnDOXXU/zHjhMY2uSA
wZ66rdywADgo9AxlVQVqV1xkxtIzFC+VaYBgdIXcBFVApobSkEx7P2yA2VonFBdfZYVRgGWCIYzr
iqYHfSaGrXVBQG3/qxa3G9pr2v+6gXkKtL8RRxGpApIHWcMpwkrB18glkFkUhlRNE/i92cAqVhGW
rzYzMLcWvo1oMsT5b8e7KvP/sifvUKnG5RPAtOWZbrDoJ1RMwRXXKPa2ZZ0+pOi9+CiMEY3Z2MWj
NUbf1bNQMQIQ/EXj3OAcjBC2ApRNlqiUod3vNn1xeWBKo3toR3/gipv7f6/wmCp5op1QiDgm6KQZ
cRetjrfXHZJLkvLqGpa1Zbe52dW6IPfUHoI6xKbKsmoM5tWsGOhskRWu1yiI01LWj7z5opdt4AQS
QgyugmUPUzfgBQtu4LSXDmELFVIHDWOstXiRnTpvsCDpfpM21xZqYE+N9opx7nU+hZx0/3vbb/WY
WECtyJZjaPWNoPLDW3uShT0mDOA5hY8IPDWKMj8Jx9WXACAXG24YU2D1sNJSoDak1YnJnvXb5KL8
ajAkNrB51DhaJLVhlJ8tcDN2kdbuXbDJuZYj9dYXN2qCjNTIMd3tnOrSyd2kKMUEU+Fh3RpZAfLM
adUvkPJBUTwMdw3ZzADy6oK7xHNzuR9yZpfq/rW6xsN7jaokDuWQR831G7lDJwnK1cWEfgijTOk+
MyYCLMiL35Fq5V5BGgpl6xN78y0SXyrwtx++uhlu6wkfEnlR3BCJ0pu6DRKgrgwLZ5F9PILBRuRF
ytS5ZVSst+HXMqPEDSdQgy2AEZloZC87ygULfV7jycEUN6ozqjFUI6w0NOt87uoIUxMx3u6pwUzn
Nmo52wQsm51Kt2G7fkenjQhfgljWZknUYOiuBGtQPRcL0r8QIG6nKA4z1Hi2oCTpvhjc0oXe/RWC
NjB38Z8/sfwQ6w/fdh+A9HgCEnMQZ9Ulf5W6JdgsCgnBKWWuSwxysm+h+6cgrysQsN+DmDaInYxl
V05hNHXH/3iVw0k9w7lUqNFUMiFV6sXBrHiVvv2xCUw5tI27O/rUt5gK9rSsYlxlZIfVvKUnTGTT
88RshDHB5iBKMekDZ5t4o0wMqxM83Q2Y4JnnQMiT0J6yL0ZCbAUcGsaQncE5D5n2B8lSVtfyt+WH
s66eSjQEdlpZTWH9sREz0dA4Ihh6EGdGYP7fD6e76wHjH+KVqh3BMsY5l/tvqzii26dPDx2xJWQ2
4MV0NUDG7ImMCyZSpdpd9UZfalH7f8i/tEwbHBXLTRUa+CGB+s0wtIbXA1pcc6v36IskQIveJF1s
/VrZeDaOuMmfuR4ntNdPdKrhSyvRpZ7O5Hp76JGPlVrJHTWgMOgw9nZHtvGNQV1c2W3e1fkaVFQM
/woDMuDF9y1Yn2L6XVLWr4K5cN9kWEkT7OnIbP8AXSabLLVDln3mxUTbdzu8sZRmT+iaq11pYCbS
IjEYF8ioqVOR5pFkEPxz6YetGZ3gmsYcNqB/Zw6nYoJwBX3RhFWot7Im7OKjkNXZP87PPOEy4RSV
vAWgcJzPyxv1mtNxAEeLQk1tK2vQR0zNPV8LNqxQsx6dG34PlJ/8TRQInlh5x43W9zcX5Xb5TvJB
36vd6QDBHQFZDnfVyGPtgj80tG50mXqr4q1pzqdll5rqIFZpFi+uE+r8PghoBztgA4kpEkopJt8V
Q+O/ATHAPKQjhIbUi7AvflXu1l1D9QqrOy5XGfamVyyOUcUZALRyFSOXoalzQygstGNvjhvbCE12
3AZbmeJJgxCr4dmT6j+a8bKPjFeZbOIJWIEfDu+KTYIw6L0FjdWUPuIAPOeUxdU3Upp9vClGVmRm
Nkqo9PI/jumv4kxEMPilCFFtF6lBvgRlK0Mv9Xs90sJ/gqm7/Ugte5kRT4Awl8vHvShqgnQe1Ssu
yBOKmlXhI0ob64S/vKoBojRvS5PjWVZxnIO6n+Y+HcQX8GmwDCZDw6emJJz12oaxIe9dK2XiI5UG
DPwVGqNBojVtm1G5zX2G3rnqQQtqjJ8NzlLOsHjsHCCRol8jCDyAKTwfWvgViPb1DOjm6chn7lxz
n6v3sH+arT9X3RpayWm3rBdy0YHbszLBkp4/rNKI4Wy15lzDc3vZYVHaRZ6R5yWWGSOU4rZA0Ghj
O8wQ5ENzCikgiqhyv7zoo+zJq439u2HS5EHZ6LkzVBeubdfi4ZATKDsUR5b8nEzmx17/qFuZJgGZ
10ZHei8Y/e6xrdsKZh+NFtYjwJeTjXr3FODyfJlLuaDIb8r8fe8W2+IYNRV/+GOVt7NbLaCAUsVE
pAerEtl7ihj1Py0XEJoo3CIXJKQowLx09ys5V478ITLnkndN4SOQecwZOa/3c9iePwD4LHiFlrCP
AKCF8gP1WFbNM0a7Tiur2DJnSicXp8sQYx58FvmtI/nWWr+4QKJzdDLEjPQc88k7JAkPoPQuGYIq
XG7EQXjKZSVMaB0BZYodMWWqZGo1CUZaE2e1l42WxiwjqU0+1MtHAddDK5MFs8+e0O+M11uIO7xs
nzmhmgCcrk8zBOxyopBeGptbYyzA8dbebu/qMTXHujSqTVPB8Xwaigv/eBMc7lhnyPr8tGYlCx0Y
iy+6su32s5jb8leY904UeRXj7XYZZlnl2+jsmYFfJ4v+elcVgMTKsIvuLD33oTvL0SsTNlgQn/lU
ya2GpntikvFtmHHB4ZNKkIfc/I2M8hxaDmmK++ODG7RpxK3/Xhk62pDaND4Fea9XnRQvKzlb5dkA
BUCWtnfLzNGu4lrfojYOKv0QCVWwwiIY6t92oVWLm8NxmagPu90gwbFgkbSL+7wtrRn7oNmjpm2K
UQk34duf4ZdGTummq53atdtx9GZ2sMXSXIgmi5mUuk3/X52u+h/7cO+wjqP36WJXCmZ7mViUnqBm
sqSelmXDvVeMkWyfSgZAo2uDqqnNmqGUaedxSIRJInmC6Ye98+i2pJm1ZO03l47pMA9Tw+veKpYI
4P8dNF8BKB5RUDipJXT+EBwODXRBK+yiNe4B7p4nxCOKv5wHgFLUvlDA4nwjaqsE/FeSGe4ZVf0k
LVSGnZAR2hFt4JcJLnu//OA4SjRessH59KPLOHqdLzPZnQ0aPCMv30IfyNTBh8yg3LZpIBckj7FS
ZB88AWwNuMB7dxCuTtM2dMwwY5IzvG/CmVkTRfzfjh/pZCqt8RZ6uUX3ol9C/m7OPfn3ulyO7tw8
9XCaPU+gfSumMhFjoP0d3q5CFMhR7Yyc/PUj2LuKW9SyDwuGnHFl/Q1Rr+ZeqIhUW0Y2s+AE3uV8
RMnccV08d1Saf5cRRi/1tx6wPerUVVzDROsaENmUNMropWylXsuBpNDcWIYfQvu2znxth+fqlRGj
yC2ZR7n1p8fHJmlXcOo7MtjYl266VhEQ82Ah4GDPhwUIkEF/NemC/WvouaBOFgQhW5Qt7XiFhlLJ
lypq6YXSvPyopmgOHhNAELFKUxkqQob6QP5VY4ES9OME5zg2cYoXtfpuUoLvPcXI7HvIsSY8901o
uNm63F0h6HTHTzRMvlJTy2iE8oobZbPYRvy+xK1fFQ3q7OoPZkovW27VNdI9z80gEvLTVyCaQiRi
oiAtCL+RCWgEjoXbi3PBsshnHfcbrLBa2Zy9qx4kn1sB1B9xqnluOlHwnYx49vg1Zg7EK3q+XUKe
OjZmqdeZ3K9eOVMp+t1sT+uo1HO5BkD1Ol/2bD4RXSNCY0SaDPl7ZZtu2Id674wZurNDAcZAjBtd
1wgqAwERQ71oWCAXB6kBWE53f1Im48zMna6RugRZ4VMSJS3U9HNcE0QqAwJoFBmVQCvN5jPr09Py
Tmwx4ToJUeZeP41C4vCjeEkfL/6fqHboXTov/DCm3xIC/UhPvs5jllYZw9q7R6CQoxgIrJkmjhDN
nAxzmxHqvCyZsQPJcsaLv4ESZhLHI0dHooUYoG82e69A/6hZomizEp0ScwWMKcaNYU29A3Syd7Pw
UEAixLDGPdZyPJuhIsZIARQ6hxEo9mFJjxPxNeAlr3BRAG8GWg6JMVR9PQY9xjn3fV5fDMPyAeI0
B1p6MwGlZpmWjBHLrg4ZqG0MAyEk1pM/bzAuq3MyUrzFUAxcKpSWDchBzuL2g6ySCg7d7k5b9G78
ajDMqsSxSTEIoHII34MZSRKEEnbJ2bamR8KgKBb23rj0xHzAdKt7paRqloq1YsWrFeiSNZNWgbv2
cYp14Dsu0OQQV2QoU/TAycF6x27e4ST5CYJEtuvmgHwG/bkCoG87MMKZfuCH/L8bU8zBEfPgkqkp
6pcDHXdAcpdXLYzD8bLvaWxZbi1ULJWpd5UTQiwADJdwWo/LlVMfE+BtCALJ+Wwh7IUVNEI/cbFL
V7oqlxkBRNg7qR2mBocD6JQmCpCHbry8bAjY5Gsto0ANzbqfvmEmMzACWpQiV8ZZafF1QUOaL3Kg
d3z7QTYF22EGnocon8ayfyl1cm2ccTdPWClbUX5moWkh2uIc7iy/bjEWhZ04f3MccazUFGizqXKn
xv7XC1jDb5CTEUkXdORsFGzcKeNQja4In7Oj0AvdMgXJGNyeX/qsMNwLAQ+X0iqQWOBFK3s9bt4N
QV28QjEfPf++CaPNXtnu1uqlEb3wP3LbKQBPilxmW+I2lsPqwOost5oKkENzWETKqYH0Si0OLCye
Lwus/zPkTD++dyAweY3vnJEr+qK9JTvL9M/TiQWxXLOEvK6EHXxJ22B10VXTOx9gL+Q+LTnczjuy
qtzEOPO8acU3Cztf228r9WoH+R3gaN5ikQAaje/hcYCyLKwZPIVM/eA4MYqEDhnykGGavBBmkwZ5
3WYtdVciXyu4o46aOtupzijxzMeTyOiqZlh/4/HUIN4WblKFGKN4AIMspjXQmlQ8K/B+wqjkmKyw
Kfw6sK1iHhixOx5un61JSnUwzbQ/7b26fUHs5AZTKsK/2DPrzFfM9CrXmNYUrJf/lLOxGH42zJzP
2aaAarkPjq+nNI205tJZaP7+xKWUJ9t4qDjSLtjlw+fiTxCvJs6Flpf+/LLv37s/Q5xE6deokyxJ
xR4CVXyYaF1OfGQ8v7/5tGDtHL7AOy+RSDlBd04Ts7sCcktBqIgMA1o+uZ8TAeo8xP7ilJYMjMNM
h8YU9hl5VVyyJJnAUTr3YLi6B/4ZPlEw7oPG4KyraarJpXCLa9OU/bVBW/MeMsEQ82ACb5O5TZCm
yGSGbYl6ithllxnaVum6EinbvLHYLLOVVP5NCERa9qbPljtGRzQ879hcZkyjqitsiIW9To6JHiVu
6F07tMijK/mAfpbBxgzSI7ZoGZFyVjLw/sszwkYwDXCjQurUwnxKzL2ZCTnn4NCNV6jJGkcXid9x
1XnUUEFQTEQLLKnSJysc6whe8ra8GdZVgZD9C7W1Yjx9t2J6i0vbG+kuU2eJFzYVQj+sA099Gong
Yh/if4z39E1+6GCr9sA7IHmgS1Q7cGs6YxVDnXAaixu5bxw9dM21iaIef7NKZRYWWZ75sJ5bsn/r
DHJl6BRYUjV1g3EYdJUCyACbAmFNolab0jHZWU0yoEBr09ureCSrMGjqA/UUfe+ha5oZEl5mCIfU
fSsnPjs219YAgj1k23MO0sNmavwQRsy7TMHJotE/d7zxFJGvKVKtv/XnL95pPxZk73uE7ziMMu43
2Ae4iEvtBnxsgvjNf2cv2OXmRQOyyPefWPMmUysy/mxJgZMYdI1yAATIMwY2txNIp/ahogGi4FJX
Bv27QcXbS1qPXg2XGO73MUOyy1+hDR773YMyXTsUadTsj+UKT4gSXOmbl0f3RMu7RCfQC21mAcm1
wmaA/yQbyyE6OOFfCF4rfl/sQ+UFkrZ6B4bGEUwBHkhmQfyNVYlo3QkeAltagRt1G7E1Rmlbhnx/
Ehe5IlOq0qImWEegGYOVVgt6NZe7es8wSN1s/TUa9ICAl7BICjRHTDb0EVmJE8LuHCh3kYh8fejM
x7iE8SWTab5g0uu2zZes4VkdpMPFTruk9ARIX7/DhhK7GbO86yY7yonWLSv3C8blAJlojEGgoINC
Q7eJ7OlFAKmsKxb4iey5d8J54X7FqEI6wyJI+aoA3i5Xo1C9UgkSO6U84CdZN2++02dBxHrvJ2DV
TBntQfZniVP1+FFJ5RDsHFD4+L0W9HpVu7C+2o794+ae+H5eD9j0aJ1MmdyWGSwcE7d30K3HjGy/
J7vFQPSUDd7ckBQFxcEiokI8w1fCulDpqvX1LpeoGRFbbTFZNE4D3nzQ+ZbXrfwS0b2myN1IncUD
J4rs/J2ApO+PT2a8MtOeUJCsmLGjXyjzLV4X2F2If6YMUfSysAq2jt6HdR/98w92Xeb2TavWtWWU
kQw8DnkkeZ/kkRCOxtD2eQUAUQObDQghd1M1ZJ+I67+VCjSSvVUonlJ6ECQZlt/6hAhNY7dp158I
zWVdIY9eCqZxTeKl1m6tgLtP1CWZpeDWduTPG18I+9PVqxEbR413drOYGu7oGvHMm2bBZh6opZUW
NopBb9LQrZ2Eq9ibBCJ5RhqtmvlwD5gSkc44zb1UDDlRTZveiTrayBTdhnBPRpb6jSndDmQBNU50
b3pEj9a15rvQU36181cNA/i3ihl3Nu6bLEYXTrW5EnEdGFBBCN6DsvHvZNvIzx89jX4l2hRqUYKJ
66JTAdoqWNH3yicLvoNdlnqIa1sqlMQMLLG+T1zzbpiKsFR5PrbuUcaJSE2mz1IjjeHjqk4mOPWC
2oMSrYrsQ/jzUh6Jndfzc1JtUuJNYOTaRm3L862fYDLHco5dQXIXZUlp9CaZmRFT0eaH72yRm9uV
YTAjJpUgMyXz1d24N3bQdi2DOzq+kk2VBkWPZpkg5eSmKrC3hff/apjYYrbL3boL59bDuoceYA6s
3rPjilPGx8B65aGHuhL+GejkOt9SsqYcttkvP8VhdS5d+drNSIH8dMJKFsoK7pb2ypWp3ir4TxFm
EDhaNPw4vOMVj8qAugOG/nQZHxAfWIU1xAWCMuUrwPZX7Ai+stdt23XRFXY+dH0vR9ZHhIVuZTlr
dEbiyPoNoUer3tHrtCOJp11w8GM3YYF6ynM5CSUPTUiS7zcwkLvIxCSSEmlwNvPt+ICYZePSaG9N
l/X2sJcPel3LeCRDc8XrzpM9VPEZLfFzrqhMZP+lv/Y2jgC2ycme0ANRBjFCJTl1+WaHgE+01MP4
BoBfYBlKCeFaP9tCuwi4WtWxt0VUdo93pborf/BTmuJyO61QBcqFP45jHOgik9ZV1fY0nSksDMW9
H0wplnWt18wmbwNhhdwGkAKT0JdSugVxIkQF2lyBdL4CL8VRV2ixkpUl2j5D7klldffTTettSooo
JkqynA2XOkL+/oQYoyH3Du03KRi5YZYbF8fL7GuRnXTJrVlgSJ3pZ4fpq1pVwT5siTtkf5J3SYf9
rtC91UFYHKSpnwSUFIOa+an6r/2M56AwqpqilIGx/ypMnzzzFjmUmKJ7VGQd5bX6SwmSC0ypX6QF
mKEwtL0jAtQeo1Cbgwjy2LU1SrVpa1dGdx5Jsm9OG8Kg8FX2EEyCUCqpSSgKDyvUDJTkM9ChRL+D
kxXGB3ZNgv8UYjli8KvSHYacye0EZB7M+XYEQkLwzAywoCVpQtmBAheDy7PHXemfvUnzALbtcrMV
OFq/6jyO+Sfykx9ASkEIszkTAwk0q9Wmmeq37EZkFOJt1fmZnN7yiPJtWgH37DIi+Lgs8zXYoUBO
eSRNiYZYh1TJMHpDVT2aem6GYBd5RVp/xnib41uEsb0Pz0AFGQ05MGoylJfADqwErv9tim5/quyZ
kdToG1dp54dumgqGGkq4znNvJwCJ9REUI0+T6AjDhkhbnqlIUVTLZMcCAlvkLQJKLH88l8uHFpGM
yuI3PLGwJErxWU4YCC2RXkSFRYCaFfDLlUI5iLUZii+j5aYL8ca1EldJzTZa+mDaT3gfefABEN4r
7H6MzWqUZ/tQ5YWIE4Vsk/qgEYClfjZydYAHlKkq0bpqJZuHHV+rY2jYCGe7eq/4yej+eFokfxH0
0THjkLpGSQZ9Gq+8Ci0vUHcQ+TDqOrf+Q9DpOBmRVlljzKAOADN7VuXYJTpGPkm0dv/2VbMOIVD/
BCNT1hj9xS/FxPMzKnCEnSbqjN4yXzGcz9Hn1X3nVTKZlUViHfPlaoV0SsGIJywAFPZ95qnjeQop
pnR9T7E/p98NKePuhSa/IZF17eibzhSLyAlMC33uVfSCG1BJ2yatVyKCWuRk0SJ1uazGOri9RqHE
TJ6yyesHTjm5NER+GpVZah8QYZ8BYnkKV/Ek0rym5cLQ5ZNjvfGjdI6T9AHfyItGKwmi21htbvMg
pQ57s0J9aUyACfqfI4PmUtUsdhuJydBF50gNS453tS0iNp6yKGLg3Yh2A9DxBBaj63/EI7q8fqTe
jC/Cm1z5R+lN+kYKW4ReyPucVA9xmSk9c4j8w2TlCrCB+8NAXr+pTPMfL/LgdZV4U4t6YSgLa2bw
7HcTIJaE+G8j/XN24NI2TG5vJeg2FrdGqF6Jobcmq0qkrM2Yf2Aefj4+i1TykosgphZuBkWAoXA0
hVa1osnIVoWEJgFnjtgBoVIxJIBHcKu55yRy9SHpZCU0JwF8tfaqH77LnVwCrNZnPEP8Xsh8PaDV
OcXsV92TeSve2/T7iQDnzcXmNdkFHfb6eEDnSxAlh0ka74D1Rc0z6sGDzeKbX+VM3iZFi+awpTN0
42b8a/GYG4JQgbKMD+Y2pfWdS0AL5K0rrTcqyQxrFpiX2U/Q99KoH4MO9/r/hrjuwK4LBh/x6loP
ckkxQ/hk1W5tYmlJKA3+eKxDYGp8v067MxpkXKrFaTdZ5/ldpCj+qt7yLq9ts02c8ys6rekGJe29
Gfv6ycXtjEhQbPbnEydrWZi7ErKRqx7eM/CCpF5B8O2PnZAePhnSBNpxietFkh1Pg+doM5y/XmIx
6SrJnP6KoEOtRDTXlXrUI6as/hUZ2RlemRA4rh6Ft3fjRX+c5UgIkk1GEA84Y1WYajLs1T1qVLRi
w4KKLsIhQany3UydqzMRMItAp/RuWfj1uobE9ceUCSaDiKPAPTa5KkrF1R50SjI2t6MZBynleI73
NHclvsLStehY1j5Hh1UKbufuDlAV7CvBRtkUbL2yyX/9s0ZN5nk4wgbZ8AMeKKCHVX7RBwYLOyIp
6JrnlMo4R0YeskzEtPV3vMDruwsMSJ0Ld8hKy0LunzetV/v0AFrkEgPTZSzGQy89XCjrtcSqfq+t
3crpS3Rha06zzdWCrLcAIx2J8bR0fq4HgvBakkVjHsG6Djb0kdcMR/qnioPxtJpEeF24CQwZMOS5
9D6IdCsxcqflYyQS74/eQiCbloq3WrlIgorHFjQrFOsxT2bd1XW9Jd3gXOR5+P5AY3jl+gzMvTTX
s/CsGX20yQn28ldhr/w4/+uM37JeMXIfSfRZbsa5NzCbffo2vkWjDXAxBCv2xmub+HQTqJa3yoLM
Zj2/AN5bZiXM75mJIASQ+DyLe7zx6MDwoHcVOULbn89x/2zAvDwLEI1JeXY4FKM8IoQFXnkE3/3H
GnlRYIs/DxMZYYmmwHqdkKLQ3J2h+n6JCpqWZpvUGzhsAgaHSGvn5+9QHrNOH4Jz5PkiYjuXVHjG
p9EygU8GKZSyyuD+pbRYvz7msvJ2LEJR0AxO0yOj5bj80DHWgiNq0/GJSjdexKYsr/8+PduC+jL/
FC5HUwakWlRbnrzYEJEXAdEZi4eQ7CYol14PEfMSfRkTSP/vnHW87TZ90EwfOIlWZlQyqz7OOzIF
0hfeIqUEw2RKbIdVky+WgrPkngJiN7WCmwdJqT6MnFLqNWYre2ZpyR1WrHIZo4U97FRwHdNcfwgr
P+9NK1yg2na3RdxKrTCLCdp6tAzkYXVBeCSaxILz5oWb5vHbRWYMbmcCRt0jbwf8BssRFmGHqIWT
cS/TIIxd7uuOe3N0HJVJhgzjcWprgWo9ePub0fxnyW/VR/ZPN5bs+B71k+QcJCmke/6szABdqheb
SE7F6k8fPY2lCikV20O71LlT/dzXAndfeJJfKM4kEvY370Eq2C2kUJHWv3eHFlOzkZkbJI06O/xt
giDdugvzSfCBR5b6Xz4eoNokjoOIILL+Tl14kEZ4MpscuXRZ0tB8Wnzt8TxITSTYWHeA0zq/yxEt
MV/ekQTo3R6Vv5TkVP2GTnkJ/WcJ5abAzSvH/uGlDacIEuz+bR3c2yw6tRupR+Wsg/ZWEQ8Bbt1/
R0AWCfWygboprYYcoCrSIY1iGabLyHlQG4o4u34LF8LorF8/2mScpoxUl+N5aTsLMi9Alk1OeEzH
UJtqIS6eUqy0Xwdk8C7PhRge1IPxgwZJOKUuOzEwS030qUtrashgi7nUDhzs1vLw7NZz25fmTxRo
Wj11SnD0V9ivhWMCwYu9H1SgLYcuySlPVvtUsDVr+1WDEHJlTfk83HOwFjCudnJ53JW3AZd1BNlm
xBmR+b6cn1W/xf+SBnyJdlXxkBqqYiibN61b1WBTaj2qguGrHUfS6KyP3qtDSPEYMCnrIlRLfp0p
KomST/6ZrJjaDz+7+pVmsxW9qlS7Ul5vyZ1j8/ao2XyRSaunT7UQFDQ2qcwL/iwYm+BKx5jnY5Em
5s59nShoMq8Tfzyxsp4eqVC5iXrSKp61PQky5fHh1mFNcA2I4jVjLy0wPQtog0vVmWR7MPdERC5J
0Hi8eRkk6Tjp3gTeYnVhR8a/FhnBOeHHokEHgv7puK9anC0q514f0EN1X2gN5lBgXqs3q62aGIMJ
gB5cggtKzgLERNQ88sinq2d1ImB0n56mB8O07xOYxTtcYtQyyLWhAFfkdfS3dUdyils85JfntQ7u
KHVUsPx/P2gxRSqy+eh4Bk+jL8oBNBRfN+S8HBMojK5qp4nQ+j21vRrcrMezO7HwQRRAXsYtfKMV
SMMohopKDqsg5RCB9UVlJSwgtkqckHJ/DcoWGoprSt+pGhCVnvpmarShDURsiTIeL2dLidXAlP4y
LOwTTFFKSh78vn9Ujl/rjMgsZ9TQG++omQz2KH4LjAIJP6SeG1lQwckeei0uQyydMHBJUAAKKFYt
erAPfRUD9gZLajDyB/9rvDv2G3u+bdFeaXy+DGRJWh+9aQI6vaYW31zUu818aM/TObS9RanL6Dw8
onZUvSkxNlxt5wGClfcwk2A3yrN2H0muPoVoYU6hHnLaDZqUirW8A4u1/HwclJhPwkcHFkp2TTXI
973GBfNP7A5fT+54T8KKmcRgZEjRx+c1chd8wwUDxlVlQ0ROefBfCN1h1Alo0jf0fHOFC+agy91y
iH/1xVN3lbExBB1avt3yLsacP+8ZMxvjNQT5mREb+vNR+nY4CPfl+xev+wwDoqtKsrQS9pSedZcz
6TaKUoNNZl1MV29Lqh0d3RMtWyWEotOdv+KasO6T08k0TlZ0mmNjZEcpz6c1eYh3JJ+EF6sp3Pz7
xE268xPVmK7BJ2KXN6EtiqcK6CB2+GWK8qqbh3P57cupX4ev1Lz64HhlPVFT7S51Ru6aQHgliwAZ
v6MZFLHj/ddyT+aYIAPiwZaOOYATZxYAHxhDcrXLfGKN4ecVQhQSLIO0WGfA+y4M/oOL31/tr9LV
Mg+TwG7Blg7dC62qz2/ueVQV+dGqf7YxOfIlIsNchYpiDwflW2A3b2c8rthSAD1AmDCPCuHpBnex
6MgvshSsnXBStryZ0LBu/SMT5J03oiL2MWcFjUqyOc9P1dqDQSD8vpCl3QslPnNmeRRaFDQTLxJP
QEsfNelDb7KyeAS7TSn2NUUZzx8lpr/r9oZEjOAhZvOVuRTRHtbzu4bJPm2W+f31EVf9U289rpJB
ptCpWn6N8h6dPayz8QBhzP6mQLJdjLo+NQGt0XXIIy9azeHhVDb6k859PLVA8lrvPcnIM8uTy7iD
QAQ7KHyFgWmRRLf6b53hLwcRRlY62w5XWxhxHg9QbgFgumA2fyMJ1yuOL7TM6lQClHv/dL6aJVO3
BPNI6dhacrzqS253G9Ggz4s2Us8DkiRRXkfEV0sXBQqn+0kGi5VybaZLKy/o9Huny3IiuXxlu8l0
fxph+3PhlIjUMIjEl3CGgVU7bnSCu/XdxovZw6N6ZbOfdS+Spq9BCq+a4VudoCF2IAlNv2mI5N5B
bVYD+fKnywnO8ket7nLRUja9b+axV3NPr+CoiEo461g8sSQEyDtp9+t76LFi1d0NTGs2wCCb/KMn
khioQTR7bzSb4n1nNYZZKMErmvhkE8gaCNoB43HnqUIvxQlbK1AY2V13fH7N/KefT5bxkYWZ/qob
n2XTbTAhaaOXIXxW/usA1da8bdk3GMaEeDt3+B04k8QPVmLFEyLExDeAJAs0VWPZII0f3QPtXtVL
nqQ3Wfe3fJ9pgnrLxP+5ZmbNWXrEZ7QJVdiVgNbqiL+76K8hI+b8ok/olZcHvliNbaHWdSYP905M
Q0IiA3uXnq6NltYu5WX9TFR2cMVUKMwcFzIvay4JB6sca6uYd9vo8WULHVX4Ocneoil7V5DXyDCm
rYqjNEMZjTv/TqAuY2hFozEdD0l80sZGP7CfcpVWQWsOz0hHpk+TSK1L5pDWw0O/4kajzPdz3Yct
VxowFF3XiIonqwoxLTs8q3COsXEZ/QoK3ycwpDYkZFMf1DllTizbJVei94wnrd1j0vOPm1m5a482
Qe9JlGVJrnL4AsaplHoBz7TnmmF+H4i2IPfwqta8zIoYST2XtRNA61nFMTezwq+/0XYqY9L0tK4X
KpZwtIJFq4BpjUiQINlwqRI1SlilA+6l9LNTJpVDpDCge/QQxrAwOjtWb0iNMnoX6JwNWYfw3uh9
ePKuVptkivkYNNgrA/SZitzx65j362GYPYzFlzrfiyZEzn+gplMraUDcT2GxqHjS4Ci0EjJfl80R
Bk6alLmF7+QgGi8Fnp7mFWSZ+2qDq42wdVUj6Qj70BAgJhmog8Ce7O0n//YVhL2aI3zy3Jk9LiCJ
d/VryfHAY9kzvmYN80yc8KI9Rr+zDd1EsRMn5mUlC04rFHZNBIghljyFdfQth73Jm+EXfR1Sz3pz
UmI5hclHJhPeqfU1GBAo76Wh/CJIOFbhv13AllmKiyT/yJJTdmKqIRTBD3tC4XpdtlWSP9YCmD1t
KZO7NhgE+yW/ykq2RtBwxjDc120OSFadxOGMr1KaJQ3E+Zz5anzuqecGo2yfD5aJOrPBifQeRStp
QcUlS7ZBhsg3k0Qhu/aOLHQ9JRpJgGfFnKTRzpUyEt/TrkRAxMVAIUMv1lj+TSpt4GsiLSJ9bUa5
Vk2aVR7LibTPWUJnnXjWzTmE7fav7BJcGr84pd0bQBNVG7BhYOYGls+c4/vKeJsiMLzHclAqkRL5
U4ucOsr/aKSTkHk30SL/rBogHccoG07V6AqQ1XTxV6TwXEZc0x98EWaYjEu+ClE9li2nuAnFNxcm
2CN+WhwF8O8o6XxnrYn6VesHeU87E6EW9SZFhXN44fdkK5Je5tPsDK9pefxzF+V8rhk/GK9ix29P
k4oExkWR8k3sihvZnbU+7OBBGMHJh3v+tgYnf1cYqX8RTGwwlf8iQVoJmMSxM+IH0qMyoP0CecK8
f/Il0o6Y2gFhyWBr5zuKHtTxYaytnMyGJEMuUkXGFy9tObAcgHlTpw45OaJoO18FNucimEXYvv7h
iSI2gu3YIjpCG2PDNOqP0QvgI5HVdSfQhPou95UjErGNbbfPoaAjNLUcMWN8SLWbU5AUFsf3vrY/
5RxdNHm32QirurkKcHSs0JTRrfsMLu5tgUFpDM3VEI7V3JJUwCrwXaq0TF+pB0+UTwb5XlG7LCS5
zK06iFqaP82CsOiCZlDeUMbZpAZY4ia7OsiUxWVqrviueYpR/H75LMSZ/Iaw00g2tjgNl0r9XGgi
hPdFa95k9Z0eO7fte0jvCcTe/f559tqosSpLoepgXslA8NCnJdMj/vfjHePT55P/nNrurcferF+r
CYEvrXY55Pz3js5VczAQXHGyi1ar8/WNvStEM9t2b6LQqb/wnv+Zv1OO6IIFWshQt8uhc9vGRGa6
OaUBvZhI3iAWOGq12kMCwxiD/j5RxOOd0+XBSzYy6fRFsmv0LFDZI89l1maxNLsvl7yHTgqtd5Nd
AoEAmnEx/HS43wlnsqIy8Jyes+smZqmw/pqB2VYz90/kyr0Sl4xUGtpORCOd6XqsyQD3vGOZneOO
txhT1QTmHxiRPPU43rJw7oVF9SHQ/4bX0R739W/1d3ZbctbQqIWJe2F3AdvquT1KoyaNcaRhDTb7
MtGEEXtmuBzQbu0eRoF9ohgV7uVtKmC1Uo1bo5a4UXA4VWSqwjrTsf31UMQFbdjdSisbr4SHlVG5
k36utz9yy4qrDlgdbQpLGMr0+YaZ0YWJpt0nxHEd+dxzBO/n7hSY40tMl5zo71k0rBaA1mbJDi2e
03qMRDNryE6CEWpuSHxfR6ZYlsfBQP7SUp9I1odO55l7O9U6TatWRGU7aPeZkX4R0i6yhU1+TdH0
H1qy7RHnRLUjfoPBDJiSS+svJuCLeanSjcvrJNW7F4NEXYLT5AHFr9wYkWYMPr+zEwyn3lreRfuv
k4G8eMfzT0CDgozwd+1oj0D57zgwSoJi9LJgQr8xJi+na1MzEQA5XJqPuGi1vy30/PP1LfMkHPXG
ayC2ZwUMQabkQY93tphJq/mlpHbPXK8pPLxyeFUt1bF9txTv0M5R9+itpIL0Z5zIGfPXjXYjjfTX
3RcozI9XMZgx2r9kpzWt69Wpkm9czK36ByWjfjtKSesZ0WUsg9w433NbODkI05s+87V7YrgUpoD1
Dbj5eOdR6Yh3OWu+KN6T20UZYtLnvYGpdC2qeqKkEmA9SRVVmB1y7eZlp0fsi+xPWYPxmaA9j6eT
xQdzfbb62hosOYvuq45Qe19vY8A05TxgXgGyNyCbzMkcBy5V3Ze2P+iUTb3fVyhzPJ71RZzcxwhx
s2AnYQYltcUzBL+712OFzcJUSvBbK/g/Kvpe27w8LfEEouy0NuIJzq6JOX6WPJGKMfNeyQASV1to
PeqOrLC8VYF+7paKHnHySNhY1NxgvS81k+egW5Z6l/smK3jWDOgzQ99z2YbhxaxkEiT4nrRwqRVR
q0MQ24+AJnmoUr4rYxdt7qvG4UwuyzVehiA1fwl+oSNmTDXsUbb5TxoTdTwP5F2h6Kk0nxz3vhba
poazxGraxZAkc6hZnYRZabtNNMJvTo7JH903ZvR0BSg+P5kOe2zxc580+ZlT38qYMbj8QNq0/ERB
YYxDJ8/xS2QOZxs4JRXXS41b2uFoqz9/RP/79sOMHQvNZN1Vkz1v96+nP7CbvR7VrYPoTAone0Su
aePqUtRbA52NjTH93Z/UikW09/fvVzgaaFqs+mza/vhlmxszSeQl8rCt/KGDJKbXGBLqY6xx/Tgy
PGbZA74CR9CIKdAzocptnfOrTvsuaAlwRUkppb8ouPrnc84yvnpK9Pk4N/nPaqXwVRuJTza8/67r
OQBtowvEwxWN+XBIkpl0d+HkavezmE6aQoXh0t+YwQmwQphqy7V59a2w+W4hZYhxGSg9VRDSXgAs
7lh0Pwo3mkQ+iwX4zCWaaXe93M4t03evd44M85FKraBM8ERRmzB+xxzwwftmSQMzV14BZpz9xanY
gIkZoRWe3YFYVZQ/mlSVaEBMPX8Cm6SLCBIaZ/j5RI1rlRa1d4MI+SoOoOG/T6OYV5zqnfDFdYAi
7CAtNZGf/Xz1Pxj3hIKUH0zK0Z2RkwXHKeVwdAxLkh7ge64k34WE9YZ+RJsyXgduBFNdNz9LB2yU
nMc6p5zX4r8Ogg0Qz53rRm2R4HuSyg1R3VYIuFAgwZ+7uICPbi3bGq47HjNqwFA5V0IFh9S71bLV
QSucpr8/TM7vOEV7S0IWXdR9F5Y97G/+LrFEWn0AsdjGFCdUY5dpgNJPXSww5fkrWOMjDLt9tINe
vo2U/AaaO1NEK9K1tIkYfy2AaaLJNwiptNInA+495a2V5Jmjw9o7yJA0Ex6+s71xInta2F0AyvwX
lF4a9sXnW618MkhDi6JmPUfV9s7qEnMB0ZFnVeA9XDaiurl947k2sZwkylMUaLpLsfwLlCbUaqAX
m1MiHQRQzcJTGsAkte7fsPNlmpIYfq87d6mO6SexMHK+38HG0+t/ieLGIL5h5BkVcz0njEhirYx/
BDLDbHzMI/ibTDHbYnF0awwV+cWRs0jNAg+E2EJ0iOh7N7GISJWGjy03MOMEkSibDl39d4FBQBB9
DEdEDQtuQ1Op1KHSBq2LHLHPuhhPpQVoRcX3UrGDIPmeb6oFAd+AAHIcgL+jPCJvSJX8Gm8iNtTM
bV6GRX18d+GiqrRpH3/wCjVXROqi+4Ksg77o7xqSmhZ1poVTU58s9PdJkSeM5d+DqaqigzCTN66S
E2nEsGgwaZBiqjA7hVhJgm+dBGjb3rACh0hvXp14V3haRl2Slb2Oqxr/r+hTa3816MaMrUjdU7Se
tWu9DixpIbnDgLnxZSdWE5GkNXHMExYwmgKHar0EmNhr34GfpV7W8t3bNPuMvuGGzhjnnfMFBH6C
i9WtRmG2Rsq1o0Hx8TmFZ3jKzK0U1jILSZC2hjMx0Tt0glYmQ4/0c7g2gjS3rYgvDvfLtzTGEQPm
SSEIJ7RA5UCjQgqpoT/njbmVTypNhyI5cj9w40J/ePjDMQnSYP95ecOB4lSU7Ur7F2wdLBtqF120
DxpzZ3hVBBZiVn1qia1nRB+o8AqDIayJ4Ec7hZeotVYDUvaaROsn/fOZKEfJqtJOdvFaqA26Yfe+
wOuZImQhm3RKyHD97uX+h2SVfkThkzXagXZe6mSTbJ2kHsiuQGQSIOSOahNx+zZcu3jDFY9U0yji
YRqsrUiQ/B4pHJZgaU8G2k2ou4zQ/HPTdO/uUPbEP3T/gagFJgbqcmUHN8EAfdw+630IvU4gZqyf
`protect end_protected
