`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
noPtmL9HRiDZQ93bIvkhXPff+H7D9F1L6e0B3N3DBnmYEADLC1VNI6dFdPQl2EhB/WxSUQIF6VyJ
sfx2WxcKFQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CM+dqqkI5tHPP5gx6cSZH1Ykj94LktinX3cpXN+OYx3VNEmx1obNF1TjV4Ii9lv1c71CQRiZuIic
OpOZDTh68EHSooVhoKOQULSZMMaQq1ojJJMEmD/3KWl4E2lOuUFzkNKXY0Fow0nN16DAfgjETI/h
TyOiqwavR4JQnHJ/2hY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
amfvr3IT4UgUDnCArXlIzdgHEU6Eyl5R87F45tEDn4ZVa8lCAlCAYQaqhFJpJaTeUPB5N0hXVAb6
BxNuqeu2omTJR4lBGjMf8hKLS5DP0fN6glVeVMBza/O4VwSnLl1hMRd2X/G6VULAtKMmCNw/8MfR
KgEK7xX507vb0Ovk40PH5+2hN1ZDTU1krCYV7piobBDA29HX9kXlJZmboXVyABsYjPa8y/95qo30
FjsgI1Vu90CmS0u7AR5MhdsJAcNHf7n76KGCaFcoaGd9Xv5+8wRLu1wL8yGIDuuYRGgTX7tBJUII
E1GTu0s96SRqJ5e9x4WHT2InC5HwOde9w42DSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iPma5lIHOuVpNgCj4n/92YtmrrYpeZg58iug/BD4meRT7gXq0kBwSCEsUHvjf/XDOrdCI/sLbwN7
qllw2ynmLI5CqA7q1WOrbD2ph7PrGEln56M56/DsembJMAuHKPqz50lPjs2l8flnP6OVYNPu5Y68
CCGYz2Zg0MNBYjTi7fk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M3ufPvOcuCqsT08/ySv26J1w9mppERPQBeC/KPANUy5Tyo8yhnnNX6eqSx3+EThYohK5qB0yZjhh
Ta+GvJZ0+fCwXKWmofGrDdhpBp9Rj05FXBIy75DmrRC2tenebqtCo8YC6h4qdOEv/0gJQbD0N16O
ZdFoJok3Eb/bJSY9tnqb4KKwDVLz99E+kdRwezT9yQ46ripqP5I95+4w48UEONDxvNb2Wbqq3OOk
78k8GSmp4szeZ2skcU16nqvA7VeOYuB1xIF8qE6OxzH+PK1+cE9O3tuWcL4G7YfzoZ61xcfSQ3ei
EqeSvhfL9fMG2k2QshL5TDaBLVxyONIV4x853g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60672)
`protect data_block
wGx7jc5qKTENvupnyITi1FjqEmFlLHAOFuV9YfwMuYyLmYDtOPjsN0WZQPXOXIt88EulhT5TqYp+
YELrqI105nc3+xUZV5g42X3Q2JPTMnU1Z+b0ueypluYBTqUh8QIFmKhFcfDvVdShA9LfKSdFjK6Y
vdqF3s8TZNljnRbhM6Cnivf9a3LQytaLRCX5T35vaGcZ32ZO3z2VwDqkvnoOOS23ae9LQWJ+Il0I
RJfS+PrkZyFeWKD66WjzJzjaTnxGTtO+0eapG5vGAzhv4xloQURzH48VgKYaCObV70qJ/8KwS0ol
mtuWkO/EYpoyDRYLSBHZYJ24xbkJqQgiZN2aF7IBWuDdJcG23GzKeM3uzgVsg48rWz6FnLdUdY2i
4n1i0u7OpgtVyoGK32kE1WBGHoaC1Ovq3A+2Q5agQewHEfax2rz3HkLe2yolId2Q6Pzo4PcaYIiD
6ShoJpzECcSQM5539O9WLK3GezHm/obbDP/aCjbZUvh2LA8dQwOkKJhWOVbrvI5ATcTJ5e80oyYa
dcYrkj0m7jTVbFNRmzCQZWBZOgpj9mFQlO/K3mwX9qSKCu2GdPEbnU5CJnIN4rTCFeehW4CSTehH
TH1oAymITYIcOi31RuoqGu0GJb71dr5KEN8tms15tF8Te7bNvjruRpC7309jYvLJtSF9Qgh19XeY
2ReAoZLVKq6F+bNxWhpgoEoTTHR+SnqwIFUhLCgLSJy65/GwHzUQ2FPssBicdVZcpxUBoSQ3M+8A
IMxR/HdfbxRbXwe5zHXD4miAI5tE3FPbsMmYVikfil8+MsFLUJSyv9Frybj43zcKyrv3tKTHDIEt
so2iYNNJZiZsrATTQbc8mYBzNPq1IZfaeAnFRoXuLVL7k+kVrCjvDKzDhbJGj0pcX7tzHswOCwkr
CDhF8r6qA89q+6rrxpl/XIFhGU17syq4bodzcg2eKsAC4rkZhLEfQMzQTYIZehPRTk7tBfKRZkOE
i26q4jgPG5y3CxtbmtfE8JH8kwkkbiMs3APDQANhSYRbo1DIFwZ2UDW8tzHHn7wExRd4emA71/O7
YBDWrK7dNmnyt3Qf1zmdpIwO6CHTbmucb9jDnDy0HWlATaG1X0xAy2scVg7FSn+kzDtLJXhvbSv7
4VWFqrl6nLGXj7Vr0WzrbmlmfOemc9z73GTw0qdKxP3DoozLTZK1d+9VprlEEa++FQsxzZchMjoL
NcYYZP/ig0UkV9rD602mZBv/r8JkdUbgiG9ePhxl55FfeaqrziYlE8i2w8gtiBwFKzBKDJ0ZZI3z
W3nqB3REBFaA7sk6OtmiPjIzawkDW1z6YfqRrTNSyoUumix9Svlg1/T25Iv/cP6mmgeOiOmDCE/J
kfBeED0Uzu4llWQdaBQl2uxBygRaTOA90myAzw1Y+JmTxO8IM2AbR0Fk6i4OURJmSkJ9jlvGP8a5
KbVmG+DQsDwaeY7XIL6uq8b+NYvtMry/mwgAmk7sCc0ATEJGfoaWyQtnbcoX7Ag9N4ARiLFBrHUw
ueuoCuLYupYK8D0sviVes4DDy2gfSd6k1qs4IXJdvKkAwKG0Ypx8nvU3QM/XWEeZ7tmoDxjUDOIT
OO4H3GyOJi0K8/BM54JtEuZKvWka0pVL744uOThJno77O7BIAIxv9GGukqc2yKKF85xv/vIZF6ra
vVGO6NiNVOHoVEqz1kHmfmoW5vf+ESw+nAnYxlUPYZH9LSH0TVrTnwdeN58EBXGIV5ZxqYc6Nx9d
Gb2Rk3IKww9lrtiyBx6hXAQka3KpY8h2DD921ieJV1eeqqv4CVx7xf+Mn7sUb8n6XUTSfZojst3T
j8Am406QAvigubADTjY5IFG5OsiWGO7BieqsgObT+4JmbUpfzGhgmj20Vx1wc6z31cAu/pav1VJL
bRO8i+orfKvPJv0wtJ+Zi8thcC2X+XALQ5kF3SqWi9H8NUwiqBSWPhobXsoy0wNz8sy0ihJb4wI0
TbbcP7nL1CQrT3zj6ge69JDRGmGbl8DvbnfxkwTuHwTBWAhQgyXKw/2izlSIOGhxcKOwSBSH8VT4
67sKfrLTiqQ4oX+in47HQLu5LfV9XHvjijk1BvGF+0wwMAxZ2WeY/01BIpOvRryh4HXNWyJAfu84
c6LpOasB1WZFyt+Fg8Z5iMX/9daOWMXvLDOHLnTr/6gtm2trDDP2ziFnf5af4XLCrgW5caP/5k3u
KtvOJ2xzUu7mPyqGjBzfyGNSTDc6QwiahmThsfezXe7bS38BQ+C3Sbmu7fG2Oka/ooFLsSsnHePE
n/xZQTp6/SCOAVjHB9H9tKe41OSj2zOXiJpOj82hvd7jJOYbrsWLhfI3VSYdUrJ9ybP+88Amfh71
nGVhQaHS/zQhuwCrvw0IsZc0pxZFmbdGU6Y6Adf6BlDTrDlCyoPZA01HIwF2ovhiUfRMu3X3MHHy
ormqIh+H6NRxNez/YMDpidXMztYQJ4NlnH3ZxPiiKv4kq9uDVLv6mn++k+Kekzs/QG9uieQdS16G
B5CxGlsW5KZcfAT8+HpYsUw7kAiVNMAkaLyE4AfXJxjsDypyLMHgqUNqCISbTe73cPgBPWi+tsXn
mbjo4B4niUa5EE9kGr2UG3o+ok58CotEEgZ3FVCD96Jzw3p7HounTxEEQVIvLdhKPlnLnE7A59ar
G5f7MUsMGEYJyqatHX7GLMkJPA7UQQlS9rMYNbugpM8cYlPF3M2UBIsE0rLpf6NiwRWBX4m0qqwd
mAxy4ZAbCHchzvS+nCpeepV7dgVN18TCjCMtbfTp1AkWVlVyVWnHKiREjZU1ujnDArkXRg1lUPEd
j9E3xKt4+FPcqw++CDlwcIrBRt3u4U5N20nLWwaQ3wn7oO2m2Cwwj0syFxgeBGXFKpgnu67+r3K3
Ify71ibAAVeAarOFVm6vaGBxbvseze6MMnCezLq+VZFVRKaYmR8y3ZFKlsozr8XSkDzM5FJehMd3
p9KPVGSDaXImFm4pv7CTxP2ftJB5DooV3bIAxLBM/gNgSoa/Ec32gbqQs9qFnGC6c8Pye9QHu9Rs
H6fUpy0u6KnKHCHYEo4nkT7WLW6zSo0GuY8dIhcfdE5ds52VOqXghdk6cW+z0nYQenQZZbGrS84x
/7vPd950cE8OpU0UW5lSEhLu/4GjfeHh14kVzihjpWB2/bBO4zL9W7wGrd1MEEYkEzdT88Wm5XGV
XgJeDcwZnfasGuMOvWzNYoju18LjvdoBn6i3hjWKikdAfsuNmQuNqOab4AFldnZgKohI7zf0hWjh
X45bXU3t62DTAxPqRh+7BwFDg9/BzFewCGZpQ353P+Ne/5/e00ShLrHzxof98b2AzmOaraNFjmO8
fthBsiCRTtTqWt6G4FaB0iW7lmJoVU1wArBNwwD6L00mRlLc6kCPvERjewi9rAFusT6zIc/irJGK
9etijfFQ2f0OjWOf0gTg6rIeIBMOnWAQf+20WVXQ4xVfSmBgw1z1495HhNSkFHvBwEEws1KKbzQx
qHqe1oEg7h8U+vzH8XsXkTAebcQTthX2UUUvntngU1kDpvfkRJwIeY74h4tkfIOGioO8+FATVgBs
xh2OKB4yjFqhO1NbfcvlT02HNVLKB2YDle2kSTm+rXixpSvcou1/HXd/X65kwrMW9GNk+RInowSD
TqSaO2GNEcHoGB95RxNyftJQRNlWGFqr+sgvKTnAbiUTM3MwRUfck1DYtm8WW6kZI3BWJ/hOQa/D
330RU/K8CTS7fHp0VFo+QhMVrq4aB8tBIX9kX98TiLokj2LWBW01GywRuKP+tR566+7xM4ywDopB
wyEP0HWqdtqiubXt9BXXJPsZpbranTpPtH2MhqJt9/iXtEnr7v+9EBBTFp7FQLw/P42VzzO7ubcL
pb2jiX13xrYxavEneqilITLNj5m7wQrPTY4ZvtyQXoKYMaN89yd1SSe5ORGfuxxKoUbee62mxHdg
NfiGCgnhIigOJdpmVtFQQyv4Mj0lPYevdox/W/vLO74pYoaqXuHYtfoF0aK7OunAfv1GbfGL6V3h
UTp/VwQTZJXZiWh/43qhEl+NttbuqvdsOT43NlmX+LmvSqiBdmGUvWp3sj/K1jxDRz9XFfWtLT9h
NsxRDlvnpvxEEjNaRNRt8z8yZuo0qiZy1TLwusnTfMsqielwpeqQFzza33pk62bWc+WEYJFdI9Kq
5oORd80f7bouwsQ1cg7VrsIUl9cf1UhVBeDNbUBVTZhXikCFEY16AsvSh8nlzSi+tmaCIGbEJPGp
EDgX9soan60H90YPEcVkbLv/Ut6AUUyBCMQTk49qODfGnJHa9ZRdVjqfyfwgnQeJaz8+cvVpg1jE
fn5MsLCsYkfLmyaMxbc1XxYGQkxTNbHQ/kDquKY1zlChKTLdm1h/2If11iXXQ2AXZ+gHb1AnN6rB
fR+SyAfqC2zI8eHpS3eSx6fxf/HcI7OciGuLfjXkDo9ak6/j5VmjkVoCuTZkvGAZJgJKicxAe++b
TKC65o0cVk/2dt3C1cJeUvxhOILCwOx+5cn2OSegS4yh9lU2/5XMGprnh63rfKThiSlPvQXv1wBa
hN4DQtClYQHDIoiHT4Ft5GQqcNT4R/RTIkMS/VgHyiCkxV76u6+DX9mE5J8PioAUYJNJKyfRHf/H
CteIIr/abnw0NUPxQufBIPsueAsFNR14NW9eqtAqwUTgfXhnOV5UUBrNacFazkvBbA7U0aIFuwnd
JZp3GhiQIF89LNZU2TovQqPMbEjJDW2vBM0MZobmrKuP9XDhyEznMcoq3jWNsBeHFmb34ReFY7xL
cqx8Qdea1F4JqqvGvhrd0D8DblaAHXA1XlWYRyVhvhkp8jpWT/GT9kkYtHmJaCTkjMLTbc+UAWyr
3GE8auNR3gQfU9fKtlDnPoCOQlXCKxUDtAFhEBNPFOLtFcZzlS1zm08fMyqZ+EI5vdiBRPvOx+el
dKZARu+f1P2QrE8LNyBv3F0JVmJW2xCGNIJLA2Ni4mVPIGKqZsVXPYhKS9vFL95yXudhxn9ZiBDD
bsI2xAn4glwYD7AvfMHP1oHlGGLRzjFGVHWvobZkGgeZnZqB3kezBs65/BMmxannnk1ELQ4JQ3Q+
kyHoJAyjRxPuZiyVpJXxrUy+mE2vp/UGU/Iyx8ZUEkkHzfB+NNX2+zwc40J598hyg5FML1mvdo/v
TtPR6RClvH/WHW384IcQoKvWbc/6chE+2jBQuT6zhqbBdClhx0joOponE92chfNTbtZB6iHf9pf3
npWnA+XeOzXE2Rrh4bqzNQFFesofTx2Z79SENA5X6OCWFLDADdzv7oC1qgVx+SixXktBhREWD5hq
Bs3dzdt+bXGGvEti17KugJ0yOep5Vw6ItdY0l27mLzIzjY1rhdVpQH2/zNUT5qzHrLISXjKx7nRb
71beNNR7e07gEHCKVIivFx9FU4f6UtEEmbAQDp0/zFg7L4Ok4SfKcYXwqvTW45l8vR1HtxfsRDOc
OmXIpk4LrHROeJ64M0Wk8OmWNeOm7CkGRgbxhP1X6kuTC1vx0/MEFFq13s3MeuFTCAUMKodyOvUr
NqSZXb1AcKG58gWIOcmha7pbVlN5U5If1oxVzZAR3xaONFNj5zXZZA85dhqberON/dnavvyQFuNI
1rseq++zxX8ak+eDnGCwvFSu31xsjDSiF85aCoRP8pZ56fdOD11sYHld/3q1GPorlGkml8XGwOvf
VJfws3/G0FXy69PYk27P7ovfs7cW0PhYfuqM99kUP+v8v8Ji6wP8fNr7crrVZlvW4ot2cTC8rfmg
pkeBCmzPMyCU5wTiLC6zpiGL0AoIbTlqdqPjPBQzpw7MNUFdwT1EhE6QhADt6jyQV3vmOoj3jYwi
AMW9pwdS4hnRbHk+WM0KKkSLcE2iyW/IIirhJwLh49uJ1G7MCJzpcmWuHGn87AGmKknZYcGqhmoE
4y1Z1pur29MyMUZygVt+30qJPGQcqFfTcTfU/W4cAssYeLo77TT76uGYrBVv1nd/vZ++k/9lYxZF
YgecgmhQhSJ6J1Wof5WQ7KIDaGxA3/j9SkKPSdaypCis8DrxE+Rb81f12F8qtupvMd0t393bKOgP
oKaL1L2XCKrIk8NU3QCP8W+kDGIydyBL7GU6n9J1FyDIyjwJP3kwYcOtFY0hMHilp06hVGnhb7md
2F2bHMebstCbSeu6WW8xXteeJhj7ld2QBVLVNaFYP9mMGSHZewbLIjBs9kFtG0sVkrcVQepDPhVL
RdD4RswUDxCNfq4mADQVb3ajajUKN1rNeQ9RCqKod+X2H/5YxdaNGHi5j77019N3qXNk1zP8K4Tu
ojcBfoAZHl09AdNvFdNWyXjsckfRQ5D5aWDnOvj5qY3covG8XCq8NGgBceouQw9cNyvxlpJoM8uf
Aywo+DjvKwS1WhRCCVnKGNPY32HMDADOD7om6p2hjlQiC5rJQZueV5ZO2EVUEMkpFx4RBwxx0SUg
tOLWzTb+bnwBTvGt01+GijsX2d1flnRotL+Mn1oNRCZlfFx7QYBAt6KBe9nVMRbMzhgTaUadhSyX
mgBFsmnBe0L3VCq4TRjQ9WwEy/F2V5XVb96thK6dA6g0jd8Ylc7h9biNRMNf6t7JjLitq9ALMm7v
ULgb6zu8as8hx7GoywFefFNmicTRBVvPFDbGFfViO2dR7Uwz2ef43BstFyEMY6Vt0riC5k/yAGG4
kkvu2qbFsNrXhTG26FanPp7bJOOqdSb6dbkqr90bxaEFI3cmzgVgYdGbbYdRBmxw0i7O0SNaLw4U
WQwDA3X9R02M8TpB3vIdUX4HZeju6HQ6D8GVkFW+8SSQp67SyQYCwEF+sv0ZBzzEuJfL8a2fS8NA
LeBFhHTbrpPWTSY6tIKjeRCP2UrY0nSVFuECF0au+P8Ney5QyOnvxzq85cFH9QU5Pyf+jRIjJarN
vcoXiGOOGclt0U2NMKl1v7ArhRZsv1nD+yASJ1nGbPaUKZTy0zBP1R4s4dsG1MdQBWuok/cRxci/
p5G+r7G69siBFIqF/7UqPPlMX2QjSzry4d66oc2Ee86yJMFjE2YO6jZwsDY+jca6pOPw+spYlm0P
P2IBpeJXuZytG5y6PZrH9PzL7NBFSliYe6dYHMW6I1yiNcYxK+wY1unHXz+VfnYqaO9TzQs40Mdo
YFhnRF0SPQVrf8V2m/s1Ig9hdn8T+i2f1XOa9TMH5qjHKMhCLBecva4nbIHctVaIDGiPihXhR59v
GWMgKpgSSzBf3lIVw+9QELg9m3p5Xff2VjPAzCigpLjfrypk/cAvufXQ9Q1eSMwkGo8j/UI6fRLk
2APRqQdUXHCQR92dGVFFMblyge9nk792dzmRrqpmEhNGIgHnXckO1nmM2xK4ecD/wD/QB5CYSJH0
de+Z9n/cNqskOOoJJ6Ha698NhaOCBeIajT7pA43xwm4k85qPfyg4bpAkt4xRHN7bFERh3OyB8ydS
cDnCoUJW8Rj28i91xIsb9RIVoxFy4R2zxwDyIBptsFFH7BBnQesD5QWw8DQbBpNgxunrdtjHro7R
NJKkwZimHk8N/fn6HUCi6zA9D9WUpZzJqhIQ3Api78U4q0Qrp8Ui6DSXJ+AgZDXx8vL9m3scrUKh
7zXaOS17rvHcrKBw+5XG4QAieJ5Lp4JiCpsC3C5BGemTCdsTfFJ7TqFGBJuM5mkI6FESVI9iek2V
uVVS0qSWZWd794HcC+n4qCsSq8gdBUZR0w0UvDXSCQhdEUlkRhst4ziV4AU3DddBCUy4U2lduQxQ
KvTpOXaPZIgU3OBW7+SN3q+ihsp4azO0ObeUc5KJIcPV70uyiNe/34xGuzlRdJMHZQUfPKdrV4QS
/5oBiX6x23+Gy0hnrRQUiAVelKJPRG3PW2kPXlb52IvwVwEGptKCnjUW0oAbu4/BdzVdSwJTQ2wY
N7cTT8JyvpAvHxTcM+HbaAe2Nynua6LEuwasM9aqpqQ9Vt6lFlJvmmOe65/1XQhcQ4zIGTiXO0km
W1+XFG9IrAKlcYWOewwSYfUxtLfvXDr6FbZZyKoFfHxDCTytAGU84y628B6QxVshJZiZGAnthPGW
dTqMKrrnriuIp8CgEGbmO0iqc6EVFt4CtMebkfUQ/WocI7OESY2irHTb45Og5gMBGZ206M1oQWG8
DXCvk4FiAPrXIztVcncrP3xs91gdFzOUTq3+cMI+YBdKfcuCU647zYq9buN85ziPDWvIYDdkALqx
SkjP9L7S/5UseeNx47CPZysTFaquS8YJR/gMgmJKjXCi7aSqfAkqX2Zi1Zm1W4pQYnCi0ztVJpOu
p+TDrliKhfXo/3bBoR0CCeEtydap3q6gn2/SOLXbudVfBnEhlyjX+2bu+IsoQGQHqGiput2cZZF4
mdFCOyJFhQw/QGL01rk5cwCTRjkgKpBSkF17uNmdWBEFCWKhbhWfKbRAkDwdMCK/858clLJpf2qV
JZln8+v9X/PtPHACW90sMDFoKBcYwXExZi+5OmVjHgBYdMxxwu5r5hl4YZgfOaropLuioPiHRQO8
qDlYPDGeEr5sT0b/QNlbCIciARyv2/4CiHCOh+EsTTJSQGJE1qtp6vR1pnW60jw/l0QXjjw9kOIr
lJqE83JCg55SeaXxl5fZe225qkVuzVDj1cIkeTPRRfK0vC005eMgo/MgSTfDzUPJBcTwagnPSJHX
hDng9qONatlpSn8xDZ24/tdRv7KgmPg9zKn42kwPEd+N3mn6FjrZ1/w+MOQ0nT/EM9h1yVOwgXeR
JM7lqZcVgvAK5/6vxzruYMRaxZ7QL+0B4YwKfSRMQ5A5f2yHuwBTvrai9RV4BFC3ecHlzo6qiznC
Lgwn/zsZtBChq0INJAnhV6Ut3buZulL7UbPCtJj5izISnucfCe36iM/WNLzQrD3IL7Ewpx6fr/AR
EFQNGQJWVoYehhjgtCXNaqCVX97yiXL8pLN+8Ek9iL96xJu3YfUKsuWpgWIckSiMiHK5gMNU/eGn
fwhkKrtWlzIox5aT9xdP2lWQ4I+fxypipvCjL8zwMerWi3mk9HhBG33DtIbzh6kCn1pv58vOxU6k
MjlY2n2eo33awel+l5qg5pD/hfzN4G+xSupnPrUbGi7jEFDg+Ck5RMtW/8ijuQ7XiAJSXhA8OoEp
fFX31wVdS7u7wjB0rOxNXn4XXTKwRLz+HVZcJ1Axd7nyERmCPgVdydZVwlNgN46WEIct67s6ULEl
6u0bcbAXXY1ixXkryiEw1hj6p7XZP6uSr79hXQ1B8PcHFnsIwWCh3I60h2pjIJbQQdtoaedKDCa7
NYHBhCp3j6JdK2BgvjZlJ/7e67zgELizgHke8KCfKey/adJhrZJmmX5GevYIfpeSsBHQPxWyOW2I
0HNLxhKDRkuKS/Q66ObD0BZ8wwQ9ZPql7rir/udgXndo3ayj7OP1t4c9iIoOREWWRexjlz0DXF0o
goTp0Z3cry02QalUn6Zd1eNJ+oTIgfCFDoLvR/yvE70x5t6i0oDn0T7+vkOFItVBhYX6SEcgsAwM
GI0wGQSEpXgqlYMRMasH6jBScrXlUvjMpUK4x8KsNLLHvExWC5op6l7Ys2AnNBmbgFbwrdlvtXxg
MFYFmCNg2jhQ9ZCqYFPnGgcxKIHwsbehknw91SeGG6FTi9ch0bXPFPZl3GpfH49Q2xz0yJs0GuA3
75kvy9uot5yqoLbNN2k2w+kLFe80w/fAmmyTbHKMcH2CTzfO4Vq2vXvW10m3ddNsZkiPuSP6zxSr
gVO0Lo3BVWxPMkfg5Ndbp0rNkBlozbe1XRPhos7qNDIbgodPWoTdfTap9AZSVLAPGh7RJObwrb1E
kmIGHyHY3ZdKiV+PwAfE7XP4MzlCk9GLcaR0VLFn7nH8yig4P7TPB3IsYQ26h6erEFuxyO4wnqwE
kSAjCOmwu9gUQDz5ca0CiDeEfpNPpsMXw/USnF+JfsuGAye+UV3D8dHoyBJBeMWANK664OQdjl2a
AnVw4AVtYABfJ20SXUAwsaHNH2nfhOR5H28BcmwPYf9NAtQ3ftPivsIuR/7t5EULwKhP/wumCl2u
fAsgWAZzOFk5ECmbcK2xXH+sT851Vyfauka7WEtjSRE5ZAO4P/R+FQenzLqjo3k0Ica70w7MPnwy
Sw4ZKv8P5l7DpwBRlAYiDCvTnWoz4WLBQW/jRxBSQdxzjlbBQQSq/ulKrY0VKrLePKNWqSP6NmO1
ZzA2I9PNaICvYjeuo5sIa+PcjoCuLYmWzjty7SfVzbVKd5J90xW39MJMFEhfGWf1g9mS27xEahSe
uXWkvJHekm+1SpoF7afMLcsz3/m2qLh2P2CoLuGNMAsbFhMkheg7/FbybhncQaWFtDiQ45ghY6xH
ACSCN+4zHPNLmnGRNtBPL8J8EvUoPJTVx8K+eik1xgqqdjvLDtSmh0KVB5tvWIeyVSpA/YgMFNx+
noJl5Lbp0nY5tHoz+Sl72TfzvbyhqWqJ9JaNr6QQZVxivGI7gWjpQRn4SPniV9p7U5fR012nVOOV
Habi5+Iyk1gLkxrsslVEOn3rHct+K4NuSYoUwYS0u9tY/VnS4CrEvPb8AV0J9FMcDtpcEKqtTwuz
DeGsZ7w5orV+ve4e4eVSy6ZtswB4O/aSXIGDZgqPJIXPYSUhMCR5tL4sGXct8EKZPX5bNAw0D4cx
50WKHI1f/57GOsWf0PZt7eCfDTsNTiDTEcLPh9Gksgu9QmhjQz3dgxGdmtQqkLBpCFTZvPvQ5kXc
4sw8PJ8Gqv+kwwg/FN2bPUTu+n+K1lvAy5IccOI3twrg5tOBUrL2RSGQJCh3db7luknAMGPW1chn
lRBERdw7NHt9Neq9GxOCihvoAQXj/Y7hXSEispCoSfjZkL9W5AM1OspsAKVCFzKbbKe4RKvE1tgg
Pc1jRjXW8qdVxG2r1xWYYGjREvhTX7fhzAekEouD5GjY2qBETvpcRCvbp66lpWxs1vwJX2SmX65J
Psia777hXgpglS4GWRal+ZIbv9i5pU8vN1kYdGRNpvRgFIh6TBnq2/kKLeZKdNACWzmN+6EGUDHF
q+sXbyxISLM5MjW24PFARUC6lFR6NUd7+fbtVnD/5BTKEBfedO6koAGr8IxO4uAZfS8veNITGICd
lk9wUdIDwFovJT/rtZXbqWFVMpR1dTGKqju8RQXOyLkKUdAIeg9DLQJnMr4r2mG49+T5lg5ImXCZ
eSpvtCU0u1w9N9hMyTEzc6zxqk5BUz7tOcRPChW4KxY27q+SuFq3qss69lOFvJVaRWRQdDd1ti99
pheN/N3La0B57PcaYh0ZdjLutMVJbV6awec/0wTtZidVMd1irwdXB8zlSh/ezkW0gNfouHGlJaTW
4PgWdSMy0P058BE8KDVBq6evVnQrdbS9tDTeCXJSaIyqZ8j8SJ5VpJ8Z3ioaXWt3d0ShReNERhnR
E5m39TDV7MiRHf14RagEjB30Art/7LXbegcrKEPGahFxaqTH+4xDU/XBsJ7vp8j8NoBv8y3Bmp5d
Di71JVjg6PF781kzCuISicsMIQz6/8U2az7xlJfiYgybL+E6WNwanekIOgHj8u9j32AgqAqIYdCC
ruGZMFLgJsSZTZwiiHLvsinQEkoJHsc5EEgbRy7ye0I4aiDh/r5Jk/+TTeelhVCsxyk3DIkXXTvY
gEj9IfZK63GgOuAjJAk7zE3fVTssXV0TzssWM9dy6QE61lwR8M5eJgXroHcx097EjbwVVFEwW+jq
/WJcvHSnIJ3pqyu1g9ONpM5Bv/Pw6zvHJpfUzHz+0oHem4a4fe+oLFjUQJaszRVDxdQZQra7/c2D
wS8ctQqBC+E4v06XWGS/Y665W7ml+ZXQb310OpiFaPtpxPhlfvSU8p8EV3Y93nbptFCjZXZFtxni
hK741tV1ob12N5AGL5NSxSKu0iTld6xCu4g2kZnkZU1loUkbY/+woGD7j89uFgyfjefzSCaOdCi8
9fGHzSAalOrtFxuNFn/F9l+AecLgHXcFQc7SLFhLOdsGkxGdWhMqPzjnhpSSZ7SLzZmE/a12OF0t
35a2jjm0izUFchuErP0UxW8GdTSAHkLK+ItbrodpCQKGmX3z9J629EM/abdX5s2Q/bItWBrMcA8o
4RRHr0oO8I+pIK04S0lHTobgtTaX5ivFQyKsZuPXaGypx04OurJTjGJmPjMkXQ/PeMGoCcZFlj6S
/9ldnv24Yu3F8Z/aiT+lcTXisIJ89TBQ/oWdeJTx8Tfo9mQadPdMZWhvu6hE8X4nDZe9KYqRyv9b
QCNd1DK5DoKW7NV5uS9cJTwqQ6Rx4q/RvoHsoovDkjijQy37x0HSprx9mNxaPdQL1NRpMBmvvrNX
FmPbUcL45tAhnhLsuTT5rJ/OhuCYJQ/iY2npxDpvxYI+tgvr97XaxPZu8kjqs7goyy0mohEa+4sq
TRGhaBxx8uDRLRPHcvHCxoW1SfLqIufVfmpRaccPS9Er20Vso3aPLf40+XM6j5Q0iLFCQHStbslB
HAPE2yaeD+kDDyq5VfT39QWh42D0Wz7Tpo/hakBsewDH2wqyLsjnqSbaI9Ok8GE/+W/BbIPvVAVs
CbUSG/yST4Jz+31dq5f4MAPfIeymHu6IZ7KMf6EosuqrHdT3DTjYmp4YCOOYUfDbBoS3vgZq4k/J
ELbg4gj8EIoE+s3yeCURfMbpxLmWXk+xf9NnccgRldnVPit/h6aUf+tDpfMvzYGQHvtlH3bSql04
ONUEAoJQ3y6u9A2G7/FrKHexnoNpyja8tTwKl01CwdWv51uEPahJEM66JUO55Q+jFC8CE13v0WFw
+Vho+EmCke34WPMWP/jscLjY5KMZphj0xlRzptLZnsQnO5uIDMtfNso+gR4wDWILsXGTAAHZRYur
QMrh/woDfAhF7QezixUNPlNpy5wMpneNhPf78adMazjI6nfIMfdbyHPCiQm65N7KJZhvkZqn8NVL
J9Mpt/FWteNkGje820/4noTxBxcFOlqHsE1fAw6p1Tqx90TEhqJaeD885x+QQa8SxpINSRkprRql
6rLLRyMnF7kRWX1aZiQJGwc/dBhVG0P6cjapw0ahlTzFzRjNfm5TL+SZQxO5USCqjydH4MqFNs8+
MQYC8twQ4mAKZTphA4vYAzjJPeavs4EOaLsmDij3xl7z0SzaVCuJcmLqITPSXUXPViryb6boG01l
3mGhpPIL2cgaYfLLPzd1te8nwO0ierjgH4ZwESXoYes5FVL3uPXYWr2DkrdMuWEUYxStq7tqFr8M
IN+YKpQJ+SxKG1A5Kg8DHYuCLfeV96djk7nS0RH0A51wLPu+Qy6e/eLFFG3yvye2XbNqLuq6cTi7
aX5UBL9MP29ljizK+PqgsYhMxt1+TQp/gykmzV00bJp9+b+kdp9SKy/KdlvZEGDZTYx0cgEJ0hgn
szQc3mDYwpoHrGSt2jhIr7cJyFZtyepCPtgqQsQRoOeSpZwCpar/UlhmAV+tmf0tCJneyI9MNRAo
JV/53YcNKZLWQc5eU7moCyb+TGZkFksuXOuv7YOb0f8cc10eQi4coTOcu3kwfRNC3Yi0X66txTdp
k/NU9z930m5t1PBl7Jy/UAtYUIot0ib5a6N3D69oIbzkaIQnzLk7jj2Lkmgr7aFl4mqx0iozgkIU
Yd2qmIZXirGV2YQqWxRWtmOd7DByeeI/yY3rfxlE09hzSgVbbzcMMKac2rExunufiyYNjrQZ+jlK
zSsmsboz0wYLqvwzT3/q9VkWqRVY6LSW1KnWUEeKnHkg+jrmxfogrXxPuwmfHMtVzvHtFpTu6rFJ
mzmwBB7mlZ16EFzvQPysXN+laCr7dMlBc56feWFQ2+A+Dy5ztvemeSBiNpoZvq60K1Kh+K1tS/En
6nfsYyrf/2EC1CoS5AYOipYLL6kUotT/aeI72OoZIkNOO0Dux2mlPcyTDe4vakiqOmB7nHeWdoBi
zqk7wUWzqiXLlxbiy3KGieBbaG/eBrfx6+ulostoc3GyIWGted8XiUSO5IX6fx0f05yOXJa1skkI
QpOOx5if2E2rbvJZLeaMqxxBDcfuRxSyzd1ICmBnq5dIYV1n4Mba+IZSaBTNhgJLdEnVwoBRJ1CX
u2/kn5+wwx8bTmuhWTc7cSCyg6d3i14pGbvI57Swkif1IQ0z8/jZRpFbszmLDUySQz10KvnEKupM
eZnOunmRQO5JGd7Xxw4cIfB0vC69C1rFRDu75x0WjkYOxLeUgJSKtKJBfak79l0wDZMa16hk3jDG
AppJd1BURsA9pmpiDfSEMMNdKHC6ttq0yWGujefVgx3Av3N+QQnmNQLzZ/GLFt/18pVsZ3xhPQSO
6GBru8Nf+g4Uy6/YvcJZUD+2k2VwAuGBpqftvEuK4lfUXQp+a52cv9teUs21Z/em0iWJ2JNyy9jQ
Z8yAPncbqWfVFaiGjvZA5yG8c460VcbXA/erYN4n41is25H8i7YNvsIekfKci5Ir2c3eBbzz9Tst
2vRdrr+w4gtFbmJ0KiiBJY8QX8pQq7w73DsC/sLP7Uz+l1cbIce9fJSsAPHnlSxOUkwQGggdt5aq
lwBlFz9qMHqTjdJRoJn4C7Z2X+rILGBt0cd/i1/3uaFa03UjAMm1JF+aSc+intvuyvC+skYaV6kX
MbwNmiE85SOkgXTgaES7yJAWNNoJbM6NggAbuvHQwja+JlSOj4LisXaOF986zebh1Es2+T+fd4X4
cdpHJAarH6ImBzCwQjvgJ3XtR6Lx2O4b6L9dtnEj0yeaO7tdCBCCNuRQ4lqIo4rAlZuZRGjypCHp
aAlYzewAOoj8Ldv3thpSwPJCKJ+ivTYe4uG99xCuAoKE012oWhktSILPV5ek0JcfcSnJ3FQkKMIv
Ui0dLWL+GHjWiLtPDRoBEG0UkYFS4BCVbL51Awez0RnSXMiwPHgZrMJS49FUfG1cC9WFOheklPL2
m8Zp07mT9XQcdBrg2N6KRIkbwWN8Zns9xF+UqObmGLccy+9ZX0SYT+TxE2Y1SVh4zKJhI4Ucie2C
8tBDW0QuGiEHdS6HLgaf5oJ3m8PpbzwpvBgW3ytnFG8iIn+MlWv7EQC7ONm4ixtDT1i60Wc97QLg
+umTzxS2slqIWu1DfE2S05cxFq9O0GtAsdqf95BtqOCTve6lsGKICmEUJYzMkOxOdTUHTwACwCXA
nXzv7HjwihPKFRu8ZxdvHJBrye2jeN26iLdTqbUMCevH58iu4+Q8OT+kI86Kpu6uIYMU2VLm74am
tVywvsW9TI4f/Ob3/bEG0HYjya/JdOkE2KcM0k+CrSy+hcYkxsl4RZ0Gv3fueO8dnR737zbhH1HV
FPAm7PyRwITfZAt8b/HkO4XZyuttsYXfXySvZuJg3opE65AcP1WfLk+o1pnv4GCAkTBbAwgLUeA4
YyjHpS6xhnKBQGjIsIG4eMVvjgId5QZF/GC/rt2Cey5eAmMo2VQzntKB1g/Sg42WGOIL7HrnmzQQ
GevaXlbZ1l8fpwZMhg8mHd2kMSQck9QVXMBgwvaCyM8ldzDYuPBY94bknI89xS7xQov4ogw2y/R0
tC1B/BgXUObrul4RH90EEh6i9XaS1A1SMKvxhCKbYzMFZz26Jl2EHZgrIdqrCiXuAXw8XnJwbzh7
rI3wL9Be0Hbh5SWpo3FU8zHA76Jpj088nAWm/U8CuKSuLPNKxv7g5LZPWc0QD1ypy9v962MgXN3F
TQVp2NIKixFP+UDjq8l+lX8+WA8RfObF5i0K2bqOBFtW8tOB9A0yIQ40yQUcKKzS3j7owGR0aGCf
8uDu13BgEPUiVQ12f+B8xOrzDWkFN5d6Ksk/fEuYhsxctO4kGaD+tQc7gsFCkwYDxV67MG/L2HF/
PXJYHuazab0fEJ7glfMa8YqPsbYtDQdZfa2Vg3U0OiO53A5tQq4uUr5VjVWwBT3B/5u2bDCoya4v
YqufkETdbCTiDEyFX3/h7OWlYRhNKMNmeqzS1QITK9PqE/OTM2TAsfTb/MlCYpCPrQlRcbdw9cbm
ogFEwB+PtmxRB+t2tr9ZQdtKxEjPPNukrxQT17d8a6UJN1HqLKQmPrTCiQeEmzzXDhheFNNIHvS1
qgDg7MQvVhlGL4XJhMMqLQ6eZ89U4N3hBIncwoynXoZCzFuwZXY/dd63KW/NPYCiOIVnl4G1iyg+
GJKGgXbRudkdAmopPTn0ZMKrY3puVuACYijvL6tZP2Ii1K2gf+E+j+6oGoepEK1Pptza0ioojzkx
gPlyvXTT078oTcWZpS2uO0Ky2cr9f8kyg+psEDTmSqIM4J104fGqjeCACeATxImwRwd+PEKgldyh
zTKOuBYUrWJ6QM8898SBs8De3Je0AvZ/pdsyUA9Z609o8GelRuX4511Vrb07BJkZx7cbB1qzqGqI
zerQDAVjVilU2digilMwXRGC4rwVi96S8lz7IpKcTVpmkfBOPcOFNP/FntGqcm3iiMdMplHPJbxS
xXpSK41cE2E5ALmJXSZ+GJH7rR11yrx3DoEcEjV6hEJ+9cnPWdN0jbFrt4tYXLsovo9X+DbgTm13
0BQJ6bgMQjEiA0hLuvoOasvEnmbgY7SmlddRvwUdLgg3gfmgs1uHm21nHgLQy/fiq8mxvoQdf6Ac
G3cjvZ2fez3zFx7RmC5yQVBMznPnzX3oeWOKxGEshSmJiyWLt4lp6Uisz67JDnubkPr38h+GG7fm
k0MMR6emZxV+bxNopDIlKpZlZhsDDYULvRE5fE9QIIrRjMzS0RGjBpg4HvU5fECU5wnJCZudl7jw
QiHzsvbxrGqGFEmMrU4lnJJoR0h729z6vj8GcFL4X4sGNO1waPcwAONJlRcLNUwMwCY7g+rEhKxT
cyDK8Q0WDochuRdqSl3J28fGU+s5ZJzkeclqB3NbXIWKxt15LugM7sFrD637l+BCBoSYipv/oTy/
zdkBmu77bsmgxDxC42e2YqZAp/5/9uqHfBW2XKRwzjvr8LrkVIPNE+sH7mUWv/nd+zkNcgL/NWwA
OvpAQZyYlfF7pLjsUnDBjD6g6ZIebvJchycC+36jpOqFOlpO7l+3cqq3Cb3q00rhE/wh+/bBsqrA
l9RJMSUP2QJFIfQSfn7zGFomuWjpgNbBRQoKY+rvpjp1g3gUiQjFK1FrC4YdcKXsSshVSM9iSkwc
QRbzvOJzDAIK216xXxVg9g8PatwSGQeeN60/ip2KXXeZ68L1VHtB1X+c+u725hjjpBQ9+RvM5Hvc
OqofBN8uhDuRrHhsNyNgueU0VLAX74tLkbWV8NvyoxaZ7kdBemK9awruhzTnqVFZC9D7gLKyOnRN
3oj6mp8NZwGZ9FGHK4+1+0On1SBcEnUX0vqOZDDF2e0cD0Aa8XM8YmfUrBGpSYm3ebGChaeuBNQ8
oeuarhEwW7cIftaFeAZK2mQO82PaCN0fWMacV83Ru5WilWtKoKO/DHxnvBFUfspvcKGkYjZpzDLr
ylRLTqzQ9AMDTT545x7Ckd+fG8iDl+0YnZLUeEn3ZIHpCU/Hg3AnU/5t17C9miNOTOBxt2318AEG
NFqz+paFuN6AI7W073jKJP9xpxSed3FixK9gNcleYFBHE+xr+PVPn8rbCqWAx/DpVyGBWBvTHEyC
5dAOb0LaQxA8yrvIjjQ7TW1GQtWPT33tMR0aaH8aDW6mBAbp/sYMcre1sjyO3mRawajzaFL2BPpM
tkhk/7yOIk105z+jvt2RKCRB8FZ5FVTmVEfNUDcofmxVK+n2Y+YhdPmExhNOh7MnCIM+eIQhLmEB
vy5dawKpOSm3u8aD3e4mTdsfQ5fz49YPN80rfz8J9D3hGJe3J6QxRJZjBliuV8WP3AOCPdPce96O
5V9262aMjx8Ah8Xs8uUqLzYfZMBk1CkSgjm4SpfCDiLeXKZEu9WZHEjctLdj5rll8R3/z138IUjZ
4PPHxRmbG4c8EhYWtpc1r4578oxS20KdrMLdZPUeZhMvXkaXut1DwZDeVV+FkZXFUwaZE5KqcfwD
cIFA9KD9B5CmPA65M5cEdO49IaEgzyT3ydzIjVw3uXe67TFUmr3XKzAzcI0pM/LoKAzBWtovoYR0
05R7YNk5FvmvBb8pv0DOhrDhlEXUClHAye+EpWX0c8AlJaYVsGZXkdP7CeoFYN7OHuPhqxiZEpAu
LgaoKIllNcAF+HEGcPoDEhlDYnOWD62h/q4NMDSRVLcoYFy0OXbln7nPgbUulNiZjWfG0IgeR2aC
vn1V7cE8mkSQKZBIxyW5mmR+Z7CaOT8+ICoBcnBjdwGVoamwGCyiQn08VRygybN9km1d7D31/MKb
Tct8qew/FDeoDuah9CFDIMkiFiyihxYPRWIQJA00aTVQ1kzf3FNneehCcb6D1SHxoauk6u7dAUaA
ivvIgaF8VqL49VBHrA+fl26fGR3/0+zCS88ZcIKEX81bSAutNfvNLWriWDN8/UcOoslICr3qTel2
kapk4k+1KF3r1hLpijf3zUTynVVF8lCaSlTPRM/+Y9K9594ESSA316mX3SfmuqL28iBiZ8pxaQg0
3UCqq7fispWJrUWHJI/NOm5KUHCwUwQ0WLl3hnK1QBRInV4Aj4Sd2s18eaeZT42aKbeirkeO+fbc
Yx2ZkW1NZIVZWHWWZL0y73GxtwS/2MW32P3OPnxmffIwHERmmc8egTPsHpOnVT5V9hyEkMlWsg1c
EluxRNtBXAujX+QR5mlGlGSpqAn5D0EaIwuWFaDYxIIob+TMoXhsiKmYvKVqKvc+mOt+dJobWjF6
vBbmjTgvRsZ0hFDOv4VoWkGOcuPjbTcn3iLt6moQFuFciQIlnjqPvVrhD8IS+05ri41B/1aNSO7X
IC3pf4ory6UaJrOEIgJUZXLZk2kyKPqQlSpDg0aohB4Zq8O9FJRHpVagf3HVC6qamA/IYHIzAp67
ABp4LtbGa671RqxyZyco5u0Xt3Rm0QtrQJz5qUi7dDithBv3UFgDxVbei/R5TuIo1SR/NRKU4fWL
7rbNf7oaPjKoDpP0NJCvd3ler+Z/1jHMs+bAkHqaDKMa9xsaVgju0kj8M0nn7wYjlDyGsKW3kYvZ
VXieyAV5l8xUOqugya2XoyvP415Swa9YRqFlOiRFG6rhxxEH9cz02cHzMl7b34JnM4UtpdYQ75i7
A5UKW+dCIUMcM8hnt0QAsnCqYnHL7bexGdB61XdydtHCXL21G37hU+LTW9oQVb0KJoPbdFGQzVoO
ppENgtrkd80i0fBqvutDcOu14IcrysUZXsNqI+A7FFBTaBEiFhsf/V4ki3vLni+c32I7dDmwKrxx
WqlDTcW9XX5a3u8Vea8bv5XFeFrz5tq7XEJORLfO4qhR/c9aimwSc5FF+xZ+coLl9PVHrrgSxm6M
bKXv+gtazdnZUDVksQA6f4Jutjz2/7lkozHI6gNTmU1kTheqg89yDNRRXvII19lyaJ11Gew5JBqW
/xUuGZfJuxgGAqRxv65lNAKbhZfc0hIXkOyZCcZvHokk9I6L/4xbKdi06p7VpL7dWboSG1emIiEj
B68lprN3CS648DUNVgunnB2U+agYsz+d49s7Yh/Ib1m1CkLIPkkbfUVLnmYR434Q0ngTmXKxl2Fh
GnnOdOo/eKISAmXYLg2lPM0XUivd17JUhZxcK416wgGbB4dAU07HXfTuBlORKC2EECmCqmC2veKV
uoRP6IYrQPl95ErHf2GMo7+z0P4xmwyR1gvWSaaJx9dwfGItGOpK+PvrU1LpajfXJzYh41skcUKF
XpMG9tbgmYrMvLFu1M5UIduKkgAOEWvDIA+o29UcfjP6357rjg12k0IBJMeW5KRn38tZMyHONegb
Cq9WF1+UcY7ZI1+dpMHWJIqx4irWVVBfbQWqSmlnQcSIKQJNe6RurheL/bLqwvpuGvkVTLs7MJ64
8oeS/fHwbGkd7vjf1qIyMGjyK1a2RtHGO2wMWa04DwMJpxYqdDaex5yfnlFSDJAwG4QDi2w4kO3A
btChoAnRdd8ce156PbmbzmLn5ypx+UAn6P3nvutsZ8qGHlV4R4wW24LNZo2gyUgaHEXUvf+ErguA
ah6VhjzL5xVUG9kzF87Kxs33khjLenzzQEiQMXUlzzoD1XGagu/B2ToMECrPsknuiL81K9YA7enL
bDssDnU/7gHPaqfolGUbzO1Lt4M/JxEUpGr0PAG2TkSjVUw8Szx09mpcYkfuOSHn3T9ptDWULQf9
k5kHFW0baDyzf2onmYPRkU3vnS6UJqNreYfCRbCTbVnSpsCHse+qtDGWg7JFIdFr7FVop2PfoCwk
q/HAxxXctyh61rPKbZ2wT/AqKoKef3iUqm7GsrWyOvyu8Ujdhn0Ld/iK38wn30rOFQU8lVzcNCUH
+MYNSzl+KO6QTE3PhzLpMc5DrW+G48w86blI0mq2Qj6zObvfU6eFnwjlijK3OyCkqZv1bE+OATqa
6+hE1X5VGL8DpUFNwqZtOVovXQMFM0d9uYZV5FSrIFD4ts6A1vYWTP6ZdIWMgUpghpnl45m3X0ls
eMCtZQWTBvEM5ngWIESwT+sv+rEW8dkVXFzsl1yPIu3mm5ZexuRsv7KaWQT/mNy4gGqLdY0VuZ/i
q7fNFeoQlP8olQFxSAMn6oNHQ6uE+COtM8QLho1o33XXGqr9uNKGlTh6+iwvnbbQYtI9N6E5+Ml8
82ED1JSD5tBVv0y6ivAsXCzExwkLvG+cjOlq81eAXeS7wiFdxQO5NlB7LXcwHDTYO6ehY3P0H3Vj
QJpuwkGo5jBvG4xUHezNmoiKHotGzFxT6LzVckoObUPk8InEt6+K/R6HeY7Lp1iC/R2nM8WoBhed
37dT2hLv6m/KNTGS/vnubLw7Ey2J1w9Aixpg7IRGnCQTqwccN6hAQQlwmP50QowxnQd+wHPm9JlL
TnfbZqxsO8l88EacTw0+5ejVxfrajy/TuhlkYDeVrGt/iIv7z/xT2zzFsKN8QyRGfRQ2Wgeaxh3a
WxbvzmAbLQjKZwHhcKr6Xzrvv2q3YNKgeV3/sjXicwkoHkhnU8ZmzpoinzG0yXc+ZwnVetS189da
QrDncLc6nJcTk/BaolGtGbMOXqoO7CSX+Shnmd/XC9ITZJ+myU+cQvL6r0jvgHVrOT8IZCYywezK
7N8ZMW/OI+ACHGPIIqG3TOYYv/u96e4sQSMN/THhRNCILLlgfVp8LQoD4ElIpjy+2HEwqvdIXrYC
QI3VxZwPw/AMN45gnRnc0xQPbQwXaxFz1FgZGdHVTKYCNJTWw02sXsMAhLS7uiElDeRA1lJd/zYM
j1IpuHfS/GJ6RGFNTXmSjSFn5rzutmoG7C0s+ccicgcjaCDXY6fC6HFxM5Gk53CMXurB+/1EfU3n
BuBcuDbG47o7e/UHnpm3W3TiJA/dCAbd2QpzI9eKWfgCQWaiMGrgxis6/AAjMlnXxiMXhe7+kZnb
X9DjxJ0mqUC+7aolaV2oiFFO0PJEvx04NF7bGkYpy5yqZhepDVtdoAhlwP2UwqcGhLiaABJzDS3E
76Fw8nKbDeMSyj9FXLR5Uj9xiZGUspQzFh4N50sBoxd46g5uz502VTdb+GZ5G99SrJFUYZUHqip6
IypmOJhRdgCIvyd1Yj9GsLM+OxnCchi3x2hBMvvp2TH086xzprgUsA2FIq6uVnemtxuyaQ1bXq58
WQ7MeNXfHPW2iZ5+0il6LnSLX+qzBS4dV8F5hiLsbdZOXsWjRlsoAz1/yvgCNu5mFGgmFVDRh1Mg
6Lz/eOtxxIMiTC82zhKBZKxHOdnjMI8mtlWL2WoSZT2Uv2ykshO3zAnpY/6l6T/r+P/f92xUPLSr
RA9ag9X6Y9AerPTR9eKEwwUNz9+GFWskDbq0ZI7xMpLCY1tEmb5N7WWc1fHqN4TZR+2TCZ5CZBZM
EIdxI1hWnwc9hTWYHzNxImygHzg1CE/RGLAmsrfba/vZk1HvY9RKGuiQefz2IVQU4rxSYmWkV40+
/IHv7pu2hht/z189WIGNDuweBLypd0WtJNiZvUBUUv8LiQOrO6CL8U4YYaBaBG2mg1XWHeJeWcha
D9rP1ZL3Zri8xIxr62hIxNZtXotBKoApnCPNb8C3yeLyyNd4R+cnt85U8vHaovHWGUMxqcXTajW9
jR/GFvj4lgHS6grQWe1M7cQ+EiGoXlthWkbDAZ0hm2b9Ho56iCZYZqtm7bLcozpHTWiAm+xUE+Xt
eYfhyxChJev7pQ8zCZi/R/pBb2luxyALIxJiO8GLlOdWVeb4zXQ0P48bJ/Scl572QFGpvjQLd7ns
z1ct6WL7VeGftWvuU67J+Ux6XPVTFGhWTsd0mvblC30aKTp+5DzExdScH8Tv3LsajJQzvHEb/TUE
MHVK0qAPwY0nEDlzdUBdrXfRdG+OZGW2F0twbRExBhylHnR5UcnoV26N0Eml2TRNx9bLgLBbnrV7
YvXguKg52tcneQIxDEtThxVIGOXAH+HDAZ3KMpqdsrnTLJ7dckZCvccFyd5vLpBvyNaaq14VMGpl
Rf88255FTHGQe1cDx9Pbz2GR9KsnI3zsa4TzVwcU/tVtxeiM+NBKSeWmsXEHBtIuvw4sB+5QdNj9
Vw9a6dueDW9XPD8ddNhTEIwqJ7RRFratN7f5gk+7zjCzzVjU7xgiYBvQcjG+PcXH4eMCeRSfwORu
l6cqIrM349tWzciBtMvxijkSvLSIGrQe3CxaKKUBQ/Ke6o0uB/gwjkwZ53WoMmd0JUC/fWHyedVl
skN8HPh4M4AvTkR5fSexyGkqTrew2zRqYygCxkd0U6ld+oWkU1sSv2y+s2kaBwwAkwU7xRoe0NWy
p7e56L/SYXsdLd/buh5soHcUc76BeArSper7K9ZYfhjrWpPVTUW6eoJlRZuDZf71gzzWHJa3car2
UXBrTsdp8QG+SNFD8lzLjPa3MVp5Fp5B58C7GdEHLha98EPizwEpnNFZhiSu/Wz2IoGRCWcLzdJJ
8Ovo2Hs8W3du1kUho0Q1Vw7xNP2X76m4OMELytWrRvGEhVG1TtNYHys2Z945zaO8F/k4tEIf+0c0
G3e3vI46B7+as3Uwc6dWhx2A+Mhge8hkCEIzri9yrY6DporKru1QkSPCvyRwIg1k5GchLFOkYrxr
0mLI5rZgerZoes1wjf3HctrV12oabhWfuIZMERq/ET0ahMikwou8CxVu4gGPRbTYLCHK0Rlv9r2d
10a+pe5lF/sQwinJw6HyDFB9ph49C4O2SBfdVmsWmLyBfjfd1e/l3ptHiyq2ukjli+5c4TyWh2BH
26DhgC/2D10S5BRH1zth+RJyObUDGEFlEJifVMbbLmavjiQ/cz8VpLnTI+dkx4ul2zB6V+JYEfd9
ak7j/xTZrUgXWAntqXFxvCfCWpOSroHTkD50kHMpwwQ8strFxSguh756m+Dk2jUg98LzudiPuSmU
Y2ZNNI3qymJuV2PfWnSHfyRFsRPgRzcKgML9jpmbl0ZGQKhHuPNThrhsyzeTAyA7PKkKCRWVIrSq
DFK1S54FNN2XTEWjqQ30fW2v4jTB89xlkTUKIrJeT0ogm/d9FF5HSlLyRp08zsFmWQ5dLjB+Mvhj
1HwFAszNajZS4ddyYvF0wzC+118MkMa/n9bU86/93Es9mzG6gw51uaB8ue/kJ6Qfy8XgAK0lbSv8
UB/Zh4+QbZWl63wXPg6MBAPsjtYd20WYUmoaYNmvmkxCEQQ3caG6aX9LiuDByxvTbynaDDaOb7dB
gPc7Nmby+RiKiqDsum/Ad4IjVhLtrEXvT/Ww0P9EAxY3m9Yzo/ddse1GdC5srrnvs03EhwHGWxTq
qpTrYxYr3d3w9asLa4SZRwMRQcpwYYo25vMIAfouAx0hAmU8b2+iU6Z289x+0uFOdkI8N5rIuBvX
+KEexPL3HUrCFgd09ikEdiiUukk0Nt2DmjvSTHZhNZC1pN65A1HrJPFzIcB98NiVKO43420zszZ8
7XWUxWgOUI4/eQz0Knyr8MiePlZ+aB7v9PFlHMXKtGbQTbH6nKWBAekmm8EzP39fbquSzRymfm2j
gaC7ZwKrimQa+b/vdIJeoQ2HjzWeFr+d+qY9XvDpHwjgAl8YyQjCRoJOIub0xBJtgiJTPueD200+
6+CMlTKTRrLhHGkVoPTnNnDPXHlO49MJd3SjesfpOzukP8e78iRxA4CRQLx3kQ8Z9c5W+SVNDWKH
pIyG0lJrIBidMDZnTjCW1KHvhIr16LTO8FA22n9WeuFREqUC9ZWRLa2nFs83vKLieItAiGt0sx7l
fbDXvc1l7n9ZIwRUgx5GpsP1SiUhEIe+dSq+YQaAO5oNuuwGsOIIKPPKcZPd7fOabix2a0RCkBld
vSdq9WyYvueeivZTzRkOgXrSlqf0B/s9sgfvBujuFCyMl8whugBGBrlW0M40e+uV3sQI+8+dv1Cs
aE/aSB46U5iVNhxkHS1y//yCgkd7G0c/ezQ3x/6FT0O10WZraTQ+SJbNAQcGONNVRYSkWoBHzpQB
evhz8G+RBbCzKKOAhUnb3CGGJFJj3+W1kQyTMLORlZJWamHjZDa4TxET8yDDY52+n+LPBsHxygio
h5o5V2mWx9SXCrsqq3egUKu+pdVOZEtrRC+ZXyL0ru0dEF7Fng+DHRTJ8p1Re5+wDNPoklJS7iL+
GCf8Y5pIdLV0XnpL5EW/o8r58fOzWrblxV6kzTSjQsHDGQxIbFvbwbjknCu6sWfvMkk0t9GRSHNu
nz3h7B+u10wFrn2EWXiMgnjuGkCVUqC6MBf4NPiPkBS1oek7DMqWqrmBJzuTQMvhMEbkJyIqRB84
0kWyxPZ51QBWAYR9tqExaN7WEuU40T9ExhzOmqd7ZZETPlXAI+i0kPZmus5lTyid1DOZkTN6PwNU
8GriOIakir65ktWORRXmAf0gbBDTCXDOTO2s7ELwSAdNNcMnQUl+Rc1jdbcusnvwccaQfNv7QC2C
p31s7fIklk8MrpIgZ0bqn7deiJvKbYywwTHM74l9CwPlHzl4iUKfNf2BrxRMwUhzk0+V5+sfPNwR
eLN9lePtFyr5iKU+FOf8HIi4vyx43P0KYbnV92z8GxbLFCttlSVS4EAYVF1mfAHrABldJP97asZo
II8QBc0NiHSjUq82zqgin8ratBCjQNwjMuWRFZNtQ+a30ly8LgcWAGHN+tq9BrXGhUZVPbf5a01l
lEpSnFjTK3kwK5aJn9wAJIaFK8Rk325wNtpUjxI+dtRoEyWvIHaPvMeEKuMQYAk45Lg8e7X9VJs4
r8Q2/fVRbF2owFDNR9cLAugqMdc1zA8qk2945hxq+vNuaZQx8OMeXlmd4I9boOc4FAIrF1zreQc0
Tj3QpeyOTANR2iVk1ui9bXbH4g76dlO2NSIx9fkzgyo0uVSE6Sty3k23sbqe2fqT2/s4ei3AViWO
fzYAiSglH1NrRB7AgRMd8UI6LkWi1mbw7fWh5+3U1Of90ETIzQF+BV5qHo8hyj+KtlkXHaG4+TrZ
HGlG58xiVAFT6TfNXc9wWdaLbggsFRzcOPVnxq+HW7Tz2cKpHI8iJ++RrgTLb76IEMabtfdQOoL2
itlF+mxHFxxbL9KWgPUMqOYYfczXczABjdmKu97eGyVdB0GvPe9NUkCw/NzQ6HfxABnEeYPsBylX
TNMrzxwNNYjeY0v5fe+dPK2Xy1586Zmg+TblL0+OoeckDVKmZa+SVbpNVrey2DcIXa3xM7pl91Ar
Jq63930GCSnWT9eNrvZKUnQh5zcKlexl3SozLEJFZmq+ZoW4xuBDbpWVFQq+RdQQerehqKiCDiZD
tu2aKhTn0ILvsCQo45s/lXPsiYFeui4KBtYcvF2xb2A0akpWClSoSK5IOzSzZC4Qi7unzwaz7bG/
C8uqGrSx+PVxpiM9FYDfQ9pnj25/RMA4FDzHawiBFAMkMuhZmkkvKv8O4sprHccUSaOCv35dDE3I
dn2Y1BaFTXS8ljp+q6fZxSbHgEir6/Yz6iWDR+pXaN1hRlLSbbASmlnohMpnHW6bdCZC7V00iKBk
W+btOV+h4KE8Z9pAOUmOkCS4PGtH5ys3RofSYtIrwzakDgPdMtY1TNPu5/t7VGtYaLHSIXi8JoAq
bHw34mvQ9DsJj3TR70a0P08mHOU4LED41rjxbcVo/hQsVZ4ssoR0aKXSQq+K/Sm7etZqvZD0JPYy
whKFCXMwp4WFEhM+GD7cAhFaxwkMExOodgUPVINqHY5fHHoReNLspX6Rpz473flez/fHn6+RQ3XH
wi8YUvC279n7F1fLkHRRjraizMktlyYuP5AsSYO68PCorSeFgN/iJb29YONNDBvn0PLjGTelZC02
RsjYYIVTAG3hd3n1bQJpYiU/5DsLFMRFRCTsZ+HsZZmk8W3ycI8ga/lHT6r+urC87mnpRzumGY8J
V9/DFA3lTddywHAximr8IHBc4A9j4msGbvwdxEBPCuDyB84CI+aZEuniKu8VuSVVKZLPFEmOR08i
BOv5qBkSRsrA10zfbsKqLtYCMlWmDmaRjET8Zk77L8XrUOEDlgDHf5bR57VA+BQ5HXQHuKc13IZy
ExMmmi/w6Mbm9qmY+akVlc85sZ8ITstv/pppnCRLMHXCqEnQ0bmRKh0P0++rSKW43YYnuiKOQn+4
eNFo6gozzFVDiXp7CwYs9jx+yX29YKUA5f4krLZnPTcV5OmwIrjdP5GokteeZejsbW7FfK8RcsIz
zwryWOouQUKiDEgFTFbJ9uqcgCy6LmBAuwbw3Pn1F3BF+KqTcuZ2OAGHzwxNY7BpBUN3KZUMmfG9
YZfBby8nYjYooH9Ay7PMIWX7qBzhiniUtVagb2nuW/+3cDZDqreK6ELS+bboTvJ46G6HpQfgVsdc
+qIcqThSvq0LVH0Qn1U+/jpN5f90+J3Q/E7piRutZNNKi8lMwifb0+F0J5yQeaLpvr1i/rhilLmy
IkyblnwsmR01R04oTOwvTahXppXLKGLwEmHiZsQG/aToEASelBGGgTj0oCIKnTBNVSL+7iMU2krc
yHQPid3HES0ULh2/nbehgwoCJPBpcvP/e+MbeoyJqsSTRiVJOWPB+KWsgfDZkaF7b1DalajqbuLY
o1npqIrVsEYy/VsYjUrFkgMpBFq3Ym3oF9xJOzJJQp6Lpa8SIgbvCKZQMHp1otFNpxeNiE9TCgLG
MRum6d+oBIeH5dv9Mf7+cG14DHBJ7BqUUCl26sgk/LoxxiJJeMZLJX85V/wfAcWzNeWs4gJVhrPV
+PStMKZF14Dd1BxU5LIMklzkXA9F+xFh5OA0JEblRzJNd2lnzM3o1AGIvbAyCQ92Gx+MAZulhV38
DmYaAhNqz0FBlxN+wTCuxrb2z872zX1w24p2x9QQypMxm1X051uoOLB6OJcNcU9i02pKQGT4Le6h
7I9CuIMeQpXjp/nK+FQnVF2lMRhBWo8aE2tk0E9EOBIf/NcC0YNdauXj9aGmAVhTpmDhdjHlTMuk
D3LKQWboHgMU/GbNy7alNOwzlbW9At2c5sFohBFD1kVadFFeTHsLB5uLhNfRaapWhDwA509vjrQf
6DaDSRTzs140mGlFIwZKuzma4val0W8Fp/LjysjPG8wdyY6Ar08fW5q+C+Lm0lbsRr+FJbF6gzqu
pFJQGSfZbl10zvpzASZkU5Sel5SXEH+X9RzL/Zn+k5fvi19U6kr/QyfjZrQaUalBOslTnfxXV/nC
r0YIkzFoYX7TQf2CGBR22bbUaQa8baopt4dyOZ5rWu3HyRbabklVYu6F84/9Ui3OiG9lYiAr6MCV
3eH5/8H1FrRg53JVRfmQxcknMThA6i+3+i8JPndizn7B/ucREGiUZsfjdZTA1JXsPG8qcHbx1eST
QdAjkCf9KqrNSPPZWQtbdc3+bZYw0GVvwxfm3FgTehnrk2ELYUk7DLmlVjmDDtGg9a6J4J+ZB7ff
TG359ixtmM+fMrd9JCgBNkR39lBGae2i0XvUgdp8z9RJU/1JNW42a6bOLRBfM3EcGpz/wl0jueFF
47imtdKjAczBLt+xHecIpXCltnWZA3oYrKXghJAluJjGso8bXvKT4UQgAl/LXpbltCM/4coTTAUR
kdSaTEkpCm+x/xzb3Ico8W0UhBi1cF/ZZNVDotvo3HUAhacFAmOhVRqzqGk/j0lb8twZa22aDN8u
diA3Etj4aIxbcTmuRRYcad3aUHIT41Mg5YJPgPjLAE7gLk8O+heDHqbb+sFxUJqRCAzL2Mf3lbyb
j9JJy4Rys/cF8uBnmSatUfJ4cfBKShXnmInmSb4deoTQGxEPt5cfVlKNhPUyyU+bPFrZKr8o4zVX
sOyOah4NZsQ0ROeCA/xFavTBLAsDUn4dPoisRoBq9rDjeefGHDlFgSUIUBKHZUW03vg1nxwZOa6x
ITJhnD0LkFvJNtg7BKzNjhvirIVpz18nYjFuJuHJfe4SHPDJ0i1L4gHl31hHOfp2CbWm+hqz2NXY
qwR+f8y4lVoWb8nai4QaqTRPor/pwxUCURuR0zCPrwCmY48+/lUYzPe19Mbyp4jtN81lPJSp79Ez
CjvckMXlEKUXodpzTDM/NeEVJd9iQ2CkX+8fZPmtkZ++2acfiLIhD1ZJJKCZ+3+IFPOkYsnuFO86
Wky0ZJI4vk6WJAwRdl/LVSjNzD7FsFsOBK7jg+iiaXNkQucKMnPVPyD445M4Qq2RQSUkL9H4AhPP
Jex51icP+aXJf5TrfnQZo8sE2UpmiGRzmtrvx0t0yxM3YNrOYQ7Tsah2AWU9OUTwJZgfB8xaCrBQ
AhFSOF4oknnT3Twvtm8suxaDvpeSDJtUYO/bzyhTQwD8HoyJAWzq524rknDjKZPh08m1VljHIykz
rT/x6Cs3PzopJnl6UPl1mATLqcq/bzTLs3sTkDAXnBPj9NyevruEIdQENzMTb4DlxhiJblf0T1uu
wlSCZnDqoJ25GHfuQerpFl1cKjROmwGdmX9nKxyLmP/rtOytyvtOLTwpcK8FOdhWPDsQ6vSHHQlM
rugYBLRFJo80OPBuuMQZEmvqAsRdxQDtFbGFjtR9t0fs0ZnTJDzu9AJQhaSiGHfuqcjIaqaSMPOa
Qr+EMBvnR6AaPsRqGJhjszmCYxwwbd/WIM5vyRxCaIFez5biNwbTVY9TusGu106sZUSenXRGS+lc
mT2fvoWWPxYdBSHncsHZOqpx5wtTB6b52iWDkEfDWqqmR9uh77LSB79vKvp7sY7XkVctoN3XEPjj
1HabmI9mL/qUUT7e95GwCdNFQd1sV02rxNarcvvwxBJtWzZ88vRSjprbc8PQtwsdNTlhDpI0puco
Bpmb9A2VP4eZ4p0i6L/KmVf3rU471DqwNgaVvO7HVfJxDQsVzgzq/jKQUkzHLxN0e2vnb+KHzvJz
shv5AHYQRIItVPkEtdFIqShi7/vPKmVilh6QdaY//ImF3ek6JD4P+Lc+wL9UgvioG0+MJ/svoJ4o
TGtEHGl9HDNpjFgN7pNBUjkLtxecxMbYxt0Ufz5YAjDLDlquX5bkwh3Sxp+YCmiyqrwiwPpK3SvR
4hamlgi3kl2GifC4CzGJBZp6IOp3vkKJdIzgh9tnpyzi0PQZBFcWRDeUAksEYm0B6UC2ILlbPr5L
ygmG6ESErUgPl/I3aIzcd7kQktJYnuNAxkDfxcZ4GoqtQ9CVyxFzgpuj1ILnDNj3lzQnAa7vPVX1
kHwf84WHjlBjdxrZPH0OGatZjXqjv8grDeFVsu/FEXhLDC5crKQzOdbFFyVKhL2RLzE4NEtI5ZUJ
jWq5a91QoEMuBzGhL47HKywtHb2LSeilLmQL1o9ojl7cxuHA2sT3Gu1V7M6NcA2n0rRQ69e6WRNU
2oC5fhNwehGseKC6NIgUviEmkcz7BWVwwWsE5+aQwLj/hMjHabDjtNQRf+7JsgcvvbsHx8K8Us5W
02iAx8edCxjqMgsL9/PG4Pjf1EywssTv5ATsPqmrgj8ydH90RLyhH3y7LllXP1xwKuEdSoKXSyow
S3olBF6nholskYsPazxwrEWWSa3BwzkzslJ7UTVtSrTtJlN3LoJ0pjiHYTSKQLcI9HcXZgNlKmnG
kttR+LcL6HdYMqfzBhIeNoh+CHWKRPMi2b6Sc4WebC8irOA62RufGMcKoUIL5VTpKvsF1tPFlXTc
apTq3xy0rWqJ/kJlvz0ZzBDR3zTLFjxvpRVIQpz05gaQNI0kKx5sbUzGR0cGrkOXWurYelpsfkLb
jjkpR77Cp5XS0aiCTWIfuWxMY5koNaFS1Hxh7O/eetDyvwv6Gw24YtV6g4OkI48ATrkYmVIbmxXG
z+n4kWqh7YKMM7H2p1kaQDiu3ANLMSYa6GhRQh3cFWMuLD98gQYWw/jEz/GBoHj2YmkZ7TRKo31V
EGPP2A+rU9XY/bDE+/KQYOSOT7zJtBjylsWClOl6l5dHwsofI908DjIMl51xveY/liWUQmtzznOI
OJ/aF1ziVTAvwqQSc5x7av+EDarpdmrjitlcSiV2cKaYmyrPVomeaTVAkSLqVnwhKZPtD19SDe4S
zAXBW7EBqByuP5gi695dmRqV5u6MhOpuY72S/8tkfAAXRAFXQ4G3XafNOp4RSfEMr1WUoNFovaP0
AlOUYLswVf9j3/bRYNQ30zXAUMKZGTkE3WL5vZwzg20mUwk9G1PUnpmEokngqurgSUqzSlr5agkP
/WXPgWjQCJ9UwAUMbKcdDd1j9ws1Z+samcuIIYwy4A4FbiGkjE9kG0jYrDVYfQnx/FCcYmr4IJ+P
8m0AzSW3RTxSRCqQsfzej0I1+ctOOWrhkxfwPJ9zIzSksXTtpiI3++FDmdiXXTFKO+/BZg4jqlg5
a+VDl4I7ToJnj1tO6ugBTvvYC6Xk5tFa+Ej30CzqVF0Jx2rqLO3zn5HAyOksPOVSCMr7QUxnUF2z
/P7skeTNXMVnPxzUCyOiSPsDzOSwUBSfDpKZXUS9fC/xN4m9PMc2PZLPXIyX9tdZ34rL4rTUsWVk
+co4ZQ2l3OxdyeHJNk8Ht7eihdQFXf6td6hrYs1VXOpZ4mdFpItKk8BvQEvuzPTFeYfj6lx4aFNn
ATQuumMKFqEbaFmKsOnvyCe5AdI68A0FwJ+OJYMj7vmpU0ivA95UAvLh/dEinu28IzbkgwYyZgJS
0B8lS1uYFTjl2ENiYN/k18cMKWK8FI25OKWkM+jY903JMflENy5GgVGpUfvEDToNxl/LZRb8mo+w
Huf1sVO2sT9Ur0JiWPy9sVuEAXDnSu+/5eBnc/m9EFL9kiBAu7A9s+BMtFgMY/oKvC0vFB0FYMhy
YetW9MY9nVHv+vXT4mUvTQSe+aKgqax6Hy4Q94sEzvHa4Gwk20Ky0LygV5GDjQgdhoBPFyXf6C3R
fLl0quRQRMVSf9x4j+RNxigmXCjsjx1C4pRZaYGIwH/1Gkl0E/rT3lfgt1U7cKkhqOYjCJBPV38u
/MSzXxHD2n1fILzjT5bfxmnJnzXW/OKALEoCb2Yt3WlKz9pjCQwpSv2ZPAqByjVGO4Wl2N3HL2T6
jujtFMGE4GDNCb+QwccPnQjaZUVFNeR2FVK+UmfsvE6Ij0Ow/nj0ZRUfPFp8i3XlzFYiiZQzhxQj
9LfB4ayDFY/Kimmsn8xdA4XcjwKeJuqQX7FJ+/uqIxjY6dkVjsDXbkiOZBiGQMiNx6Vht3/6XfZd
x4ovMO2036DW1yvhA0UsINfRA8YxBhDgPl4UA1Edl/xt9Lm08dn+LmBtDqXB2JsjkaANYEHzGaYi
dKrH+Lce1cv+2Vjncj+XwnDx1g+F0ce5EI3P2L6lQ9aw3aJki/Gd/R4x3MKqsRIfejSpMr/SjSrl
/E3nVNk2hE5ewlRpvUcaAg2S5WqNBlM3hM1yG5mwTfpOlFL12FvAC7PYqcscWL37oJksgDGP7c52
XXaLD2Ud5vpzN6Sld3WeOe/Ol1NGD8iWlc0+gK04gSxUOqnz/ZFie4oi7l/7Tacz7cqyiHhS8D5e
g3i5vpPWPHUEqELyDpvc01LIyx9PRojUavON7I7I4J1a1eYyEduX/oqoBWCyq8D1s59miPPGYfHT
4VJ+u+/GoIJbi8sSLU1ZGbS0mMx0bkGOueuANjTv7UnDnaUs65dIE3zv9SGQClJU63LV7H9H/OQl
PUDATxXO14J7fkIjykFfqxGACwsg64ZWHokx9kkDyUr8D3PpiN0gMTSEZzhKwLPSqP7adKCQdOcb
2D73KOQ+KYqBE45fFx7UKxyGbBGg8XlhLYVtKSKktYTjfEpA8HlF9lGR9+Si9dUVjZJ1xzBBiNP8
HQb6FdzMAsXtuSFO8FBD9rIBKpmo1lWXSwb6wNcFA6sXC2i2Tq8CdoU3d+xc+EpgUEcxkTjKUvBf
t3ZcVtXybTTay3lOzDojTX1mJ99k1eNd0bed5v345pPAq/MVCO/dBcgUL2ndKREIgsu6ypBi20zB
UyLjAGBpKRDBg7zLYcR80Bc+GI260m3ayZlbv0Njes7JQAx1xSUCLqqNmwUBMk9eZtOmJEvTvOIg
oDn+NKEqwosyiTshUzLLKJpVGNQSwHt6QkdxHDEQ831A978+eu4cfqZG5m6x5f19W+RVnjtoRUOz
3y7Uh2qcEi47U2rPXwQGR+AqgCwEp4jPBcIRYlGbAaP8fObMiPciuygG9MwAcIz3ke/BuywJVAKW
k9kxUWS/B7K+9sZLT+sEy9zSrwh30oyfCbZ7AmpoFaF9dc0AZafhqvx1bzIBseLHvD0I6EMx/7Rb
kQG2Bj4YSk0hsO5XzrpIfjHXXOMWwA9jB0e2WfwrqDJ3UswTgVGf/UUlyga8W+fRYArDQBC/2Fmq
tMr2aTgcfsKjboUKbls7RnC/JkLGULjjmnIK/AaAD06hUFxLQ7dWuUchoKskhGs4HmWXBuAAY/Ta
5FNmsVznNyE32VRWET9cfAS4QZb52TeD5U5M/GrLfLP66Mdi0B7NOf8y0GUN0Ne8fMtoMPQifJW0
N1lxI44nMerBdL7zEj8KpL4TwJUY66wol1NEJaLt38kuNvnUqbwytKT91Rn1KVVnicRdsQl/hqzW
ZmKYcwY6tPULFqf4vj1HTnDkwIkx4MIzCM1p3Tzuvvh/1/4wLqKpgwGiZEvYvE+UFmJVJwr4maob
vBlowejfgaCnwQTF1BwG+WRDRn3r70SMGco79ntO9zoSGPxeGFG86KEIFDNJyH3s9aPNP6UF/l/5
z7+ZS+rmd3kFD367uw7043lnDyqB11J3pi63ShfoWGFXMRRjEm173yAmpHSrdfWyVTif5NZwGwjb
xDtewm61X/p9Gsxdp/PALoCPPDWEDr/ZAfhyZGJGlJqWHEVmz90ZHZJWpeGqAfL10J4U3jAvxAr5
uHnhbC/a4z5kzBFHX+MHgTLFC34g9PNhX/8monAA1Gg2ltllD+3TYSFZ9H4SNhnWTc/FhSLW32Ny
jdzExvf44Yops8o7uprP4deWWPj+t27I0hyItzHlLEyBSHiI5udqiwVtl9H1TkI6XR8JbPAmM+jR
asVMOkTEXkLrh4ZxBECikMvfjQtxw0E3q/s1dZhA9Lk2mRBVe4Fh4qjfZabPPBPEGKN9Np6MrG4W
iow1q+yg7VDC1oNNGM1jmmhjtaSAD6X55XSkLR/J6S2cu5/jaRVJsyNEWW5ohpMwOUzxN6K2MGDL
HjFgSF6cZdaTwtpZCc3cEXK1TwBCrhGKTcNPLCi0SxFBkDrQ90mFSGHKhsMft0Rbon6pT/l1Z1wJ
+Mu4a8HNBEJ8KUt+bNkzibAsQ0LKL6StWJhiCU71DhLbSELUrLnLpObzTvMaRgE0OTg98QEgUQhJ
zoBCOUImEPR9REnUNYyzXFdB3Ha1e+X8fcTqBsuc/cELpLQeUgUT4GYeAsiVOzI7BpVfjrPBzuyU
pmXgS9AltLr2k6qP1jgpMl7h8uzGHdEZ9ZNUfQpickfp208rBwdi52Dyd8tlbSBUPPJnh3u+ZzMw
Y7Wcez+dpnDxJd5pBQ/DM2TBtoMq+D93ZdhIO3EuE55ZciLt4u0SIhC8L1HBqj6oSHJTLz/XNAq/
oA9iYZ53ec7t0mAPkAq34kJfmdKmBCtcJ179XHZzSeh1/qD+fvD5KQLBjzWXXgwRv25tUOpGPMwB
vFrYlDpCHoYJ3vVQ6F9Z0itbXGKx+kJRuIBL83yZ5jSn1ZC0zcczeAVgKrdM8uMtzakg1liIs7CV
ZD1oITFR+pJN3SI/oHmerIHtDC3RJPxvWbcwY2K3HeWb8n9t8YXeFufUgOyFd/IUoRGlkBJtZzqq
GjMOxs9ctkbnnTXFXKt88cahPPAUyqE594kOD8rWYo5DvzgeJwbtMJjwrVofzgp1R+MKFKgH50/E
N17n4bhuWmUnGp7UmIPQy1pbSWfMuso5pm3zaKMTMYB3mG4J2lenqWtjTHhm2LyuDSu3SBFWB3n2
vZKBsdjMieOHAeYtStAL/XIQZmAcAHbzBUNVq5UpWkQMzSb+33moNgYzTa/Os90t0BPPec0n5RyN
0mqhXcfEOIf+rqdflyjgnadCmHpoGMLl5iSPO8O31FRIaAj2ZFEAAAD334voR5ySi8DpwDle0h0z
rinkF01vRwjjSYbGuYJwQpz0BVOiIDQiA3t/uX1HOl6t/o0SZM/3srvBCBfLCPZtYgk4mZP7kxob
eAx0qGkWRpFBpW5iLKqCKzVleQ7VFW0aSy0nggx0Y3aziRsZF8OU2W7B9jLc7722YfFz6z5AJLA7
9Qo2kg6Uy3ZqwV5SUI7OHr/oaj46OL0iz9ieSv3NN7zxGmaCnY0de5OuBvykzz54mQdJzq5jWY11
lo+QblL/Y6zw1CZWtGdsU2lqXoUeQ4lzo8LGITqPqPPAFRKWxfUWrhTdZo6Jlaz8L9Y/BQp2d6Rj
a5I/1AGEdMMuLe2ZZb6wyIxNilYjOGPQX9Z2y5WROS/oad++NP6KIOpbXOv45OqFbrKZk6CYJHT3
kFJKmXP99u0obTOyKSMkt+WfXfBNjNPKP+ysYH9sgaeWQnlzXHgMZ2lt1odRt4pj2PiPmyfCET4I
Wr34+5B81Mr9l5EjVOwlxRdtHC397wrP6a9EjCqVuKzwTA1EZXJoSc/ZCvZMiTKf2lANMbueFR9b
qTLYjnoFHkpFmxPdzxUIPNsjyhlRLQHDGrHu3wS7+h25kkKpWD5YIXWKqK7kaBLmtoPWDj8S4Bfy
lt3hx2vfUm0zCX/nG1sZzfqRna69x1sQlHBsXWbZCz01luGwImxYuMNUsK1ztAohQjeU8x+o3d9T
ih/ZSul39FRHL+ajvUg+d3za3i26KsaADRYY4Q4J4HXnRD2jKqBx6O5zpDg/TyiPlUCOtn5uGy1y
DNGTbjYqsRa5o03pvuTrGs8uZzitGYN6mBL8BAxsiJs9WqHXhwDD15pRIx8lsTr8kTBNycbpRBdE
YbICMdeKe6RF76xsDlnT37sazIaQZXXItye+hv0htfTF2hyl384hqMZc2i/Hz//cMIOT2TnfImhx
EW2hF0zlBfhLQsTKP3qC74e+7+9TeRuEY08AYVkDhAS1sJKfKwn90kcvJ8negoALAvzs27B7lZ0/
8sojEnL46WB/yyPaxesAIrl0wTvOCKUdL0N6kY50PIjPfcOisPsOkSUXKKYKzFoSxyZWLoXJco1L
YUq76paR8jU1Fb79HNaImKRai7AJKGDMBdCxgzms0uATtjMYpWvPCkbRJ5r4AFPv9+64og7+NXv9
sQzvgS7pznBqvG97FIoI2wp+bByreMSHYLWYbhXBCYI7U5W05AFqgHB/dDaLdl3tUTkTbHtyELBc
9AH2+fYbJNma0JysbDyndYgsfAjiwVaJ8OyBg5tjJqEHypYzSxSLhKfo17IkiHbWqFBsqBIu8kSc
HYCCGKm2gDElCWgvPhGkPSpkX4wQklcfvM+8YFYPa8pBADe29c0H1rmr3nOTAG/qiw/Hy8dYPAv4
3fVwfvFsg11SWb1VMeVoX0U7/Z+d23nJeIEH+UYdW7ii0tRXzu2h3Jm2zK7ydawS+urXf5UyYsoI
ioIkUf31UyAb2xI3SWRlTXz4LzYJiMVwaAQLJIwuPzZS9opWoTd+jnt+BKytI/qbMQmJprEdO+Bo
5aQjOJ093lwYyAvAeKjLaTM6GWxzOn6evcLpLDxalkcD0tCfK7AkGHsNTyG/UKUHf9vo5kq3rFbf
TU3Qhw2j2yZPxNfnSIhEnreqn2ZRxtB+cjpfsRs1+oA58eDZg6g6kpwRROkiguTV1reeeHVmwV08
Gso8QB/xt01oL8V/D/WGnkV+eoZGYSpIn6vo1R7tHHEgxl2f9R/DE/HoJsu+viG8nmHRmG2UnznG
AiZK4AG5GIe+RDF187npVbr3auirfXf8h29v4jXtLWLzNj+YbVblbm/isUaO0pwxZz1K9WoAfEXT
UAdNIA4uykg/lBxaUkbe6aSl0GR2cMImMFNfsgZNtRe5lm30nWaD2tvkLEAeNbqaoCDamTvlSddU
PylmUh9nhJdPVWE2H6YLAB8TRRhF5xWpX1YrvFQ0Y+M/J7n7c5Bb3Qf+CDZ5kkXQ1rtpJyX0eQPS
qKyJayXyLZs+9wvnW/9CTughTmJkVXZe54ZJroLNEF1v2OdfcnSHhGfZraEpyvdcPxwmjgaDzayw
R3lMgfzbAJTfkJxiiwI8CAl+Nyy8yLuy8I8CorWmnGMEII2j7sh7BsL2Mrq3f8Rc/I1X0f4/BwGi
Nu/MDhCMVomG7XkGzYOj2najfIfJzcFQdI0gSfjTNRUCQ+XlxZxD9BukwhC5XulOZ5V9WJJqQB+a
5sm2akm13/GXL6oY8ipL8I8pHxmor2gpypkzE3mN+28P+TvOH8ctEf3gZrisKQnrTsb3b05dZrg3
O0QJUAKw4+RTdbCsKrpBOOcMUJHblV7uka0i25AsAH0C4owNepqaXcUa2xkgA1HsdEaFs5Uga0iU
et8frr+in1DZBFp3/a3lunmiLKXIWjKBZIcL2EuMcohgpIwJjVLAGjGCa9qpAC1JFE9ScrCxrkZW
eEW3EnmE0JURQx4f3lFJ3yXZXrixPEqerzU1rmVIuUPcpyRskyQEQhs9hD6Z9+bc2M4Amhca1orC
CD8Wf+IGylFxtZSMUqarpTXOVC4UlmcpNjSXqqIB5Rly+1YC+umrmgjgd+vknZuco5vXQSDKSz42
jmLzYY70vhl9wuJX54WAsv6cWrQ/yrVcmapVE+XfLPCEgftJFSJ+Gv5g9r/Ieob0XIiSCiu5F2du
AzWAAqo1RxJjAcpHJalzv6T+QI1Y4h5i91DVahYWpCEw6/PRABqF/yc6MugvKA5PbtC7VKnb9oTH
Jn6IXUR9xpObhUmLy4pgZC8EGfHkdykBrB7zjO5pBg85TeAxEh020mRZvO54a7vxwh2bMxyJ0vb0
uW2utDuYdWNv3gDSnKhXkZZBHgDsWmIZlF4XPoGi+CexOr1SoOfV5pg5AOdch4A2t4He3uP2KvR1
8VFNTbyq3d09A7YQB5W+ccjR4F2JS8R8nVeni1bvdopEPN5xX8KzRMET3BRuhF02lfqhMN4XnEgJ
fAbi9YJml6LiOr7X5WidNxK/W/WkWeWhIxA9wqfczGh9j+0NAFvcGrSL4OdJir+QIV3tfZ5p6Oqb
R6h1Gj2I7AOZgwCmo2KbyUoLkVfhYAWiI2aky6pO/cv7/X7ZChFLIXiZ02NrbT7P2fkC9855/d1T
GreCjLyb3VI+sMH8Pe5tuORpdtL3S8+Zm51yZLQM8L95E24Ye9LG7GHViyjSVpc7+VzJ71uzb/Kb
9R+ZfbWTFRzWr7dB9s7qdjZ7fF9ITVZiua499XEAksTxIBW/Yp7g08A2viR4CE/DkPllO4d2SexK
/8DXR6ADd4mSzl8HREFCWkGrwcSXZx+reAszUJrE00pzTL+srw0bQ1v1f/RMq4Fzi6EXp8yHK8Cs
FMeAVo5kQvo+y0RqXYPKvPk6H3BMdIPDFFmCVV80ihtcqY0dwAiP7z6lgVGLS0t0FdKgli/xsL3F
8xtK8nx2aotWvoJJ3W8gSmUX0Me7mB7Lz/T+VGtol3nwEaJztwAiRBdRB5X1KjqYOr+OD5BfUqgL
AnI0KCMSWtAmNYNHJt/p3WW14woYXMbWbhGtPz+A7dUaoOxG92tSo3rVUtwn8cb9MQWQNGuUJ38J
KjHluUunt/zRNcZ6tyvTda9tkqEdRpODYKHX9DxdAZ3tQrSK2OwAg/Tt/yZuS3dISuAoxtOlj/8/
scO8yVh3JftXpRueLFw0wgS96CMblSDvR3LqqCS2uTuBWqtlT54KfmrVjRm3jmQ7w1MLm2QqKVPU
3OlWU0vhRwCpZiEjzZwhLq11u1Jei12fegzz2JvrPooaXyhGZWZzUv4OIa2YWuDKA9EpNjT8uQIB
qrX4fCnsJRF8p7Lz/qoqBvoPNTy2HzBWXloAIFnAi5eHP4U824DpcduMnc03yTuPvUP7BMdNa6nh
u99rQgyiLDBW2Y4nXTHKbHCZwEsPL6dnPdFv3EycIdnY3TiwO7tE5IHyqZ9qLz+aIFtF0bbCy6RY
GD4E/vJKjSy/1ME0t/csFPnuhf4tprB1dvMpAyDn2JQ56gh1ArIIK89s91z81UfcHhkdMqSrTeyS
q96WMBInmt9cs1npAyZWjLd1BvGwl2z8vcxpZiZ3k9KNbM62jaEc3JS4RUqDJ3s2M4Lq4eeCPRJ7
URY0vUh0qnYMIzw5XIeh6XHipjeTbSx72ZlrPVDNYuWNUlarJzhfU1LJN0ucyETqHAbiOUiG79tJ
Y9JgTkqd5DruGwyZdLvwEriSXT2sG8UxPCMN2zRo4gYx12p8vj9HgGFIs/ZVQmdlaah6UPiCGxWd
8iq4GynzEHFeohE0vlmBMHQPubNrcfObjN6mXgy0Q4TY++DZ6OfzH6aonYrKjFezR8yP02hazHlq
h9vmhFkT4A0SQI61DbfIzK4EMji5athM23+dknNqTmpgnXhdVNl5vIKX/pyKGwK/TKmYla8lO4hD
VU6ecxuBcvlcPV7npFQqtweWZC0epsY1p7NkzfqutU6AFPirHwjz/l6j+gAaCEhUQ/bMIH7V9V9e
N570Nk02v6UcC0rLZnyPZvvdHorBQL+03kkYwCEuTiS07yEBjuHLMID0OXxMkUybnNvBIKDWfUFg
7bHnP2VWij9YmMLg6ZbpJL3dsTjQyGUD5y/+5//rJwtFQbb3cbzD91FeU2KM3GtVTxtNTYmL3I1A
PiUcotpDTKMA+Udw7bShzfl6q+c9AYZFC886A0v/Wkf5faVcLN29aZSl3SIu2cVT/nNKBINHCfg9
rAFTvEOKkYTN0JjtgDxw2/vyIQamKegNpbn8/m53htfrfFRC9Aejy3waaofxLO62r45MY4ykuQ1E
mnI+8ZuHPmFy/Zhm26PKh31ZMZbfrh1v26wVfoSBEflMdtqvrmrEbRf2aJ0/vwY368kvnb16njqz
ylF3iSBS1xkggYjVlpKO3j4CDYNYyseKc88ZdWHzcfcG/l02pzfAdws1siIw/kR/FRVjlR921PPP
RLa0AVu0TGjRhF+ey8K0GpIipzlYMddWclVJ3soANlLWokvoq04AKHRMEp7Ok0nXOb1omvZh38CB
uyRSlKQE8YlM9//L3VwGaDRfuTwqeas0PoPUvzc+Ak+R6YI7Ytvu1v9SdmpZJ++zLX0DzH9eihDD
wd/WT0TEzAypOINcCbJHsKSg8WKe/YKh3/bRbLnw2mGm/opmGHU5AWhwDetI/VAAfkJ1Gtd7lWxA
j8bwP7PyTqwDfb770BoVbVE61IDGe/9UnP3qGkCqyOtmBpmYmuPs8j37Kp8z2AZBUrWQJtQPu0RP
ZPhFj4/x0b++72jRS/XLLKbDRTHhdTnyBVtP9rKclSml8UBwMRgr0JA1yoGvUpYUJtn7shKQclxi
gU2DH1aTHkFkJb0SzMbRAggoh4QUrReK8Ud3aex078zxCDh+1amYiRfJBYrPtZDI+OYXtjgTT4RC
YVtfEKwGlqiY7/w+U8qE5K9fs2VVJ/qHT2D1dh2SBjDmuiKg+Q1zHQDNF73TRfJBzFj+VDZ30CER
WE9655mupYOAP4O1Msz1WEe1belqmKkoA1d48Ex05Tnp9mnHmt3x38qvs4ID3JmhIyrm7Seml/u7
9ml02qJ30DVxqTkSv372UXoxmG+N7r92mA9x9RvYtZFlCP0S28eu3Jbn/Yh5RdvMabtH19MAXQsp
TT/T+AlcCeM0xQA1M9snQL6w93i1jeAgRktqNUSj36J3XdX7NBOyO6VzkgL7el4isfx8EgHfDHPb
ILblniVx342IhmsWxs91/GBJfJjLe+DoTj/q3ZO/Yj1E6SkJfHHylGdH6gxiiORZ24AylrH7ZG2b
k9/fYC1fZOJJohmgVHHcpcCCqfB3Ukr1jTWaDumSLIT01ltFgU1q6LJ+X70qVRuElof3wvI7m+FI
PU6skXmLQdvUIot0PC25eh/d6Kqr+jayk223vEh13h9yTAAOnRcNuiQjxmfpEdIE2OjTLQWJ9Hbs
oKVBJjjf3jnkabVyV1ZqZy21h/MNrsger4Yc0NKVzxxGcg2bdTLOIKhRmneoCcDaOIfAjHzGB+6x
7KDsL+twwF16Rr3uSeOJTu2Z+JmTg5RrVzUfv6e5HmM8akeqsAGD+SqCHLPFM3/EmH8eOXiMFszh
JiHNncH737b5jdY0G6fvfiajpcUbocWDvWMeESkMiCP4CJ/NCo6f2poNNBgoyi6jMuBN3RftW9Rm
ejEc9IQ9pnnuY0/jcc2lf7R6K1Znyhh7WEVI4wpUZyKtyEAUPdsocuaLy3oAFh5pLzSvnEcuMzqD
0TjjstDDf506Uhva5R5RsYvfsco5nD2LEbV+XrFW7wn9msgapgmypbUwNmBSdpscYNAJUo1EqCBX
P+2pn1HB9tyLPROSFVTdyDDZHEbberiezmQG8IhVCcB0tuArRsSu6rbCAn2uyJVxIcUjRrKTaUnU
JBsadjwupCS2X5vI/iEkpXAOeDEQeKQ56/edboRn12V4r4gVovO7syvSggagUxSKSyJVGvUzVIof
UEr8DPCFcUr8rLZNfMI1X41iyVHzbhw/oCr50oNHkqI8VYIUvQhAA6vmS+1ANMjdakFXvROD8v7Y
q6FKFzw8EA1xrHBb7+eDs4uCniiPw/4dCazv3FlaSO+KLC75yL/tvlyFw5O1n2Ox++GqyjVf/bAu
gAjFQ5RmbWfKrn0I3KOI0Q8BTOs576KfJXrJ7XReqqxKP+IDzSlnsdQQuELnIoPPQrHFuD3N7yth
2LJrrUmaWAGBqT54pyM5tzP7N6tAj/aftTXdB9ZpzwAGYQB23KD5HIwQznc5wD1/EH7v6Uw0D/C0
Zzv5jxX6xbLFR6XO0SDh2oaRUM8xTktBINecGx4HqWtdvyzDZZHIWVyj2GhRkBjR4dB6ckj6+8Z2
3Xbwdvb5JuPbVl8GVL7Dx62Zfwq4k7G+5YN/fOJ/vv7mR4xFM6Ih688uhSKwnRsQeMLHim75njbA
0BU6II0YKfApIKfYb2clIvd7vlj+6FwbZlhoLD8fTxEsSqzk+xRXXi207b0w0bbnOA7kNuTL7wD3
GfakXKwQgAukBPJ4glTACI/wDChjFbu8fGZls0AF/L33uOp7kOzEUaiTMSE3/Sv46zWeNy24c6AM
GSnEBu/Jf59p2rRiGCwwjmFef1muzsRuZW2K0+glkXRThpbGJyMJXYxmSMETBQfg3cXih59NyiF7
MOAb0+K443mtlNTS9iq+p20vwiawJsFTyXpijrASbwyDCV+rlSSZsRTNuXK9GX1CVy1a76Y43LGU
/GwBRfl2O9/ZoEzjowz3P6gy77fvuUkK7b5OXpEPty5JRYM5YqErfS/FONL+GPVWQ+z3L63IZCKh
Rm94vd3QQIMbfYAJ5KkyX3Xvyax1mAaxH4/2b+cQl3nOJzVuD2RqMTRwAfM++pAOVXBDUJ6zOSO6
37kB5C5mw5J72MickimNxHctCkU65y4PNeiUdJvucOjKYWvVZR3FG38Jut+rpFHtC6bCOqXCZSdM
Vr7eOCrRQhF/NeBS6aCSey6KGg9AnLI678WX8CCzr4OMoP/BS1QR4Zg7x42L+C7nhvUiI6wNhf/p
QPfLTQOJFP4Q5xOmcu5MYR7jn7jxSwY8YQm/GiauiH1aCyOiGRYD45x15yTFLfetXfHgWKjCi/tn
MVbPqe4bnUXhO75cOInw+t64Ll+hUMzjxwDm//hVNZri6/klbrzffBycHp2CDHoCn3IfU+cvkMil
Nq50ICOrHC15CnhlWtmtMB7jC+dO+RYQQyL5fPd7QTyEH5oFmJcfi24zYM5aUshbPwr0lCLqWpe6
Vb7khUyJOJeaQT6ZtfZxbzWjk7iWZcW+MS2KusbibJqfoGh8p6iOR23RHsgHlhhb7k5qSMmggyK2
LiY5tB4rjaaDDORXZJlYvF637u3TFLwtUQtjpUu0YEoXpIhvIWqNOvPHN5CLKA+uYww8iQuP2mbm
mac4z8hBn01edrzHiJFU9IHyvzGibcRgp7XwDwdBjVXMwIkIul5hBHJJzmn8SCcfBdAHhqVAvUH8
RfuhCvQabOVg3WvoDc/qjOq0lXKnYKnUGemjcFQfz2LYVhHZbFWE6Kpm0qsTT9vFpMw6PQ8UV0IL
MvuXxZuJohljbALjMey2eKqwrE09hstFWT5ZT2nDCYd6MxlkxMl5ykYVtyhq93rJFgHkC/Vxdxeo
ZQ0d9NWHs/bpKsbdqhw9RJAGQjXmHqVIGYn8Sdp6BGtpWLP1dpjZJ5mOYEb9GhtGakC1ksAjh+QA
DQS5QEbRYuM3ekSj9TYAH9oQ2JkHap/RQSBj8uKUYpZ7tNqSSeXGjvOjepRR7zwpZnzOXAF8MqPg
4Hl26/pW6YtHknOIHCWXCDU5Vh4OakyNPzezm+bfu1FpvE7CPeZCWk5EZxIBMmdCwkAwNyi726y2
d635A1CxmY5H6FuO5Wgo5v8YZWG89eXPYy9VG92XgBv5Mx1z7BaPXRA+J63oPA7AHh9dxMbDi8yI
es6mcGRjHZC8BBGOzIEEZ0t4vlwZ4CjEkvP2sjvpKAfwzYdrz6ELAnKVKQ+Ua9eO45vEqHb9AXo3
SunNZKx8Zqa/Ct/CHtYdb5IFX0IP0Rvz7tyIWPHEwH6or5uWBkJPGOPXOknxwdW4oxeeixog8WNh
N7y4E3ug3mmJWZ4YWxIFyZ9ZJOEML/+s/LguSZ/sGBR7W6hGj5l6hyEW7Ed8drY2YxToYs19bgt0
vUWYqh43xr2tWgnBcHcBd5Ac3YWhOx8RYjSyJblXsWnO59y8dLXqHVm5Z00jXAZBTx7hxaKrpwNq
us296ChtbyydOWWJjU7hTO62O7V75e9RV9/76dLExFn0Q2PjWJSeaz9KiIWPurA5GE5uM87cSToF
6YCU3LKQaacqq1HIzfRB5givkjIa3/TVy5aiT+KgGTWQuvD9rKfYpdizIUAEfvpYNhaFvj2vIbi0
Dgq69sy9KbBRGW4gAvYdVo34yeh4zXJcI/+810lcQwahdolIcRoYqH2k34rl/p/sqJmYOcCQv7D5
/vu+fJFYFc+Ha/JcFPTZZ8LYkHTN36eU8h1XL4EYqm1Rh+rV9GYBauosuDpfyyZSiT7VEcxnxmI0
C4zSgYw8LbdavPOyiCB4mOmzVT2XIAYyAwnAFDJ/eJveH1PbeWDRTJ+5uwX3nXMQ89XVFSHbOs/E
P2eHji65TTRE5sPFjM3zVZdgxTnhkbtLu5XLNVGJRcdqkshUDDdOvEEiITUnFXo/kbhz1BH6BeXO
+2OAr+AxNbhb/tw10jWfvxpngrps3ezSSkRDI3NL+vE4FXWuaIN5rpXmgDPSNbMJuiLM6llzeEWY
djLQWQJ1ZcNsB7NlenL/8QTUnx68YASbaedMTPRuVyyEvO+a9s9bUwBGDEOK6zxNUHYmHoPeUGd/
FkZVEgRrQWtk5T7z63ASD4PRYumGOthJkkOIPnDdled/FNcH4OfQVX21CWfsSjCvVDyCAYdv/756
FW0zX4Faed7gI4aNTEsn/YSRaB60kDbPJO74KBX0qnrD+szfa5XfucvLCsNumCtjJIH0Q+JnD1YH
VAtPdnUI3m1U4x1DNDcVUTSAumLlTn1PBr1/t0tZNYFYMbbub28zYI0rL1bGiignPs9eqjTX4lMk
nT599WF2RmcFnYKILCv3syITLwtsR0c+9DfVF8Zjqjzwp1OSB7ZJ9KSFNOLFNp4pI6AmEckZjNUe
mdKqRHc6KTcO3+yls1UDWiL6s84NqZKN3FG0WPkG/8gcdtJjWjkLiBdXRgd0c4F7wRmke5JpfQIM
IfJEckZmlEHdOJadb/28us5Ql+paQ+D14S8a0rnC3YxNLpyiDwj+v48bmk3J4isSdmhqWUsMVTIc
41ZyxAi19mHFXWNhrWyvruNbqjQ/SheilivB4032Jetf2VqDwE/Bni9dG6HV16BLUcBK9XbBUbPG
9HzVRBFfq6JgM0FLeHc68jhEH7UCr2fdtuTArhpPctx/8CD2UKjaE0K4LpD1JH1vI8QpBiHzp+ik
RvE/pnWWdBRmnHjrMkyvyQokiuSaTbXUkc3l1EdO3G4av9bX9VECFFVOPsuRkQLOr22mHPJ7XJen
vw447eJF5PQtrdh23oRLDftrOvPMh/YjqSs/QeA8JXIt9AxfuaiEKGaDamdR8EwWhZ9DeZ5bFCnE
w6BOAojc2N8A2PaUypmPIx1hw2xDi4wNujrVHPb075DGhMBRkxODkeA/kx471FKFzy6KZ+OCPbRB
0kYxKj50bUuXcEbggcsZSoxYi3pxkd9TDQ7ampvHqZe/JWl6nxTadblpReu+6csBGGvm8u1KiNrq
KGHOO36inw6Y+8AS9HbrtSWVdbTRFwDo48OEqr66s6NZEs0OiUPHCOUUw6SFHjwgvKNiKzXN0x3w
Ekh/fVjt1WGN8sW1XDwwGEKlM8rB2MmlSYdz1KRx79Je0htPYxX3/Dk4UZJPWUwTFi1Em23wkT2y
9+7LK4EAGxsyZ+AxAb8bEZCARos2D8ECJmEwuWyZY2BjXuXmq6dd/vja+w9o5XdmNzZxhwPDX0ev
ZDjGryE7/ErKshxevJGg/ZvClGYi8Qqgl0nx3Zv3+CxewRXw1h3kuhkBgqQfT4dBO5d8yWN6g/5C
iuFgVGO+TqkOwZfRry18KE+2PYpJNPwUGoAXzIRylRYBboO0Tq4rcaF8SFsMUQs/ctoL0bZnDIzD
uG9nLalNm9/LHsVv5VDGjE+GmMitS2S/5II3fuT6oSEsqLRW9SOtSiXYfc7lgdvys/PbXrLAJA6Z
aScoNyge79L6RDLWVq41YaG8cRjkzhtgdLP9TEHV7MNher23rk084kYSAMb8dTihc5Jt17EhgpNz
WPi04wPhK1d6ZdoR6EpWfC+7S/ZJPI7mg8idhynGqHFHwqGJS0UoyFUWN6u2GzdAnEEI/IRBY8K8
vHGc2qTtYRkGxX9nbrTIcmldzgO1Fr3u38LJI38/P6gJcBV59ProxZ86iVoVIydVqNfbJb3TYfk+
OLnXcWh57IW59fT+e+wcmOeBVCX5nXEnGVi+YYB9+7X0jiwUkqZ/FEXegyaMlSxi39LATLpZJzFw
GHTgCn1yQw7DdvQsxowja+dl93oWt1XBzVylJvPnrTl1GqG15qRbjttpTw7O2GXvOIIBNrK3Rkid
DELn3erejEc1kWX1nhAwIVjSGl4SLXt3Z6BnIHtNibgCVTE4UehQ0nZDyqDk4IPNkyswehglcpKK
VMnekfpnBTm9MP1LHa9GCybVUj9hCViBAdsaHsTOuBiYDapwtdfN4nG4mmPvolFeRiNGY1B/a+R6
ikqD9LklZLx5TrULqMlMU8M9GHJdnUGCtU6dspvbkEuHw+8FCPtqiVM2861pCqOThEEtk1AWVBME
ZskafoZ6pvx0JMgSt3Odjjxak2bIoFAkWNEfc7q+5Ogi+BmDF8QMrXbpS7YVFJVtsmLdTOxQlCr5
pL3gSYvN3jvaoo/w0YDHhOuY9RPyADP90ZYGHqWoLGMTLBG6nDNDtd6DYXAFCLor9z1HVsiKiF4M
Wu2ZdJXw/s8IomRixE0tEtPlXrtjDgNokrnIJvRoVc1Jgvu5keKTo9Y0KrAxLU0VMzfa8qFJQxUc
az02xVpT7qrStBoTOZlbsXVG6ET8rroMIaQiZkuXLb82gy+Ar9FmiHMGjmb3ksgDfgcSvdNDR1+c
vO0pWuC5ZCgu+nY48O8Hi7vZFrReWbjA/QmZNmtcrXZg+OT4BgBYRUen1SdGso3beVRH0ByiCUQ6
mdo+Pnmy0bbqUxM+e5SVtRwtYFwLfEJePwia/vH7Qt7UXQWUVMcc4PD6rFNPm5IjmPPlb2UWCFNR
16cBG4sWLildB+6tnlPTCOQK2SzGrECpORPWARiiSgOK6mC9wmIi5LY6CfkV6ksStuuyLHd1SmY0
YocbY0i8do7I0N0xCqMyHY2JsIFdc0ssDsyInQGL5p6hj8ZmfumuKYGAy2xzwPyrkoD1KYTH6+Mx
GkZVCe6jjIiXBhd213HgUbSe/o5iTFxXBMtokaUKl0onlF6KXYKFRRA2isarbaXjgFTDYnF+CqG5
uzpWBYJ7b0bgKdYEPUL3/MmaPC6as4zWTLkTkH0R95p+rPSsQCOWbkylL+GRP0WzCmFwbsdQkAnk
hMPqRpL0mjm9p+LfgD3cRbEUa5AnEK5E11TuzIaT3dWgVrIlh9SA6b7XuPsBg0Q4yIrlVzfQCmmM
TiltrMvivvMNdq+1TNMIUk2ZS5/A7HewUrbrwXE2St2edbw7wIi6dCnuEddPBKGWebPQXIKqIdfr
8EPWxrHK2yhtrW84hHH8Oc6jjnHbUbTT3izmMXTWDxVXXaDn+0MoBR7zZlGWuBCQNz91vnxELDjM
Sr0XIjJnEbMVmU4B/8MttaFlrGwGGsbUV0ngsuA273OcU/z4gtBvt423oUE5+Jfu6YbcK8mEI/9Y
OyaZd7ExiWqwTaQtcRVHt2o6WZSdbpd3MpL/gcaIDo2mNVQBRcdEplVAr96IHDO8jEXHqS9hHaum
8qvRXhe75UMiz3ENVEwntvg8InyCgt2z7Ogml6BKLIOUMmoG4Gc5F9tssSOpaAHH7R5dpV4OBX98
zkwEJ7LYEZD/0DXKusvWTToqvCKJ2Sn/S0b/75SwBZ5g4pSdHKwUhJEvkx6O+FtPgLDaIW3XZox1
O7LIKLkyJqzhq2fv9s4k659wubhAcWH88Amm3JbOoIzdKjUW38R/gr/wWT/0vuAzKPnbKJ+FOF64
C9wanS4Y2Zuh4sJ6wEMD5IXeT9cvzS+eQ58qCk9npJcJgN5bVbB0Qqd8DeTjY++u+729J9aLEvWM
Rl90vJX6RjDcwnaFlTYGw1hQiO/CiaS0SCY7TUD5Rpy85e/GV9anBq1cdxGy/hXI3NG4WTbxBxy6
Ms4vpLHbOvmFN7h0HA88VBqUsWiGe1idN2dzcFZLzLRz6iQzimlyMumWS+lpvVdypzHKhwhHVRTG
sn7ySLq1GpZiMXi+i3COssYoPlf0mD3b4tPWJOJanIyHaFMDF/IUYySX4hAH04DH8e5t5hRP6Ekj
ooedIwpUJKToJ1X97XwvQse1bsD2VGwIGOs4azc34MASeL+Osbx8t2IE7VwJE3yLkeR3GI5kpnJn
S4dDEvPcQhJksujWzoDW5pldjpCEk4YLeu0aMKrcUI25g4pSSm6ubqR7EO/8NAMKDeV4fieKOmCf
DUs9eIYN+kBv0AWa80gD2micQXSpdx/wdJzILK9s0KQc89j2srIrHBmkSCSEe3Y/VkCHFrYXGNjz
kenqXiwmx1XTMgkaLjwYARQKrW7BZFfmeUG7hUp8Gvb3nqxtVyqqkc6/YhjqyBHnULrKFR0CODgl
9JAxExqu0wkd5HL/fwjforkXD3VNj0F4+3IUq3tBNqC3x5Dc6ISbS/SpqVsuxPhni2tBUfYSYEF0
VzHNFuIYPqxjxmvWbZGhKuy+TiMjrgRU+2Y20WyMt1OnA9+iny9E6pj127aFfMpXcvb1Ts0Nvrik
1wndCSlfmRm8w9b6947MaGCiswvqWyhQJCklwDrkYvOKjeTSg2ariK5IsJwJyK1Q8eJ+B8nYXTaI
sGm8QIGUv1TleUL4DY15Cejjore0i0HplGBYKP9qrTzbefjZiRXpTRChWUYNJmv5Fh/NM02NIpOF
hVMV5VQxxBbNzc+FIxcMO2MB63xInLtptCenOqQioHTj1dRrYAodAozxzApTL0wahbajlTzC/P80
kSTshvY8mT6io7ekdpFpR5OgBZA7Z9CeDwPFP5BoJL+NUR67rbSYNK8EfJMQmNMhoH0EhYRjHUQZ
sP0km94heeMhDqKAgqfdV7D3BOEECkL085v4dbmDrOFTVKw712iHq5aK006E8orbdl96CaS1hRtT
owmBiZSco/wjV/wgkmGJAB6h3txCBr7S9oun3J/zUDJL3nq/tlOY0JSEEU8vj56Xo0hAXkLaj5gA
xucMJdn3PQ8CMzNI175YvijsxfnpNLO1FWXPSrCSD+Ou3dzePElJ4SW4rvBJPM0kHlG/VtoUp03z
Jtfmlr3fk5CXzwKXZbfC1GA56uXBSbvZ+NaYK4tx6L4srgkpjnvXkIxltP2NiFEXGawYPd4zfuRl
YXObDSpLWER2xugcNiuKF16KhkssBIk9y48Kvo0o16IGeL4+oY3fyuy+QWUpexp71FqNAuwAK1sD
xlaATLmqdIgIQGZkXPgJhANmMtmWXc3/6IGYrUxSaaCnHKdVASrDw66jTe6PK/egx5yVDz0+2MB1
4uMhNbmN4VkrAV9lqNMlkFfp3hT2t5ZvK7GcK7d2SJr00yhx+xRfISNYP6t9DrlUs3pWfSkfSKpz
qK4T+LGfDQUVLjPmCXjUiXiCnYW9n5LCxW84vYdzI5FEzNLlTuNtTw0IKm9+Q4b86j3y2QtovumS
++1c6FA5chdVe3ncMqj/Tr97KHMLvpE7XupNLfm55o8dsibcRLMrbUp26Kmn+K5aVpZfMy9eaEYM
mHFuRd18TdBAh7cWKDpuZ9oTQPm1liSLP42LfL2ADJ8ICns8rBpb2NbbWgxxBDzkYk1cGfNMR/Is
DnvVKBTBXli0gMxLd89lFaPIZf7mbp1SsgD/PrM6C6B8RfQ60UYeVxjW7/FYv1dqjP/g7KhFMfBE
EZuodhgiT3VHeeE/iI8v4FBequwV/7+SwjoDS3qKtROvv1e9fVFyFCHwhgXXDhbf7gJEGmVgtBYE
oQX9v3dR2iIm6uLig9cBBsVdyBR7DkexBGdpbZfvNUph69y3bp1hUfYF5GM32ltBaoQ3/v9FpHRN
XCMmCSNlE8F0Yc+ldxdl4QxFzyaGp4BG4P2OV1X43LVxcvb4qjoVY9YxtUZMRcvg13JcVsySjM8Q
pGWihe01MfNQtogBOVpm/dtYxFJRxgdohleUnmz/bN95qLZuxcF8Br9xs2RSZtl0TYb/y+nK0mTO
g2vH0zDcYE8cTasbrai6VbckZpLsx/EwSiNPaXtttiTSEmlSuwhiYjwffObOIC0DKf9CHfs+6P9C
TKFYkbTVJP1rf18XarY4hTLKcIjQqVdnesuNQd4nyrreuxiH5y0sCF4ZTET8y/SvpfZgu8EJZRAm
ypEu8o0VyXdNRYvCRD+tvx5ZA7v7P1F5M694sZlpY4DBQAtMW/78otdVGdQv0n68d/QjV9TxCuyV
vrxXAi6N0yykBNYrhbwz5n/uJ+n4BTgZFXJfYLl1mVTKUQB/DfVIfh3Jmhw3scDP9GtptJGe0/mC
WbLUOF+N4avwtRz5Xo4TT/DS/j+3qSOLN8n76TGdZxDzoetKJxbmcqKV+rNQIPlB39f8PGAmekC6
twNsxwL24jygIKTMucolqKBuz58+I6H8UfoPds15K+MxsTOxbazb7KRShrhV0MVYyoZU7rWtpamh
Y9SRmewYWqJeb9Bh72SVhDsCeanbmbRfK2g+jcAM/cmrRFDltmysGkaxZ9+qFr7yrcursAfpKdYF
GbYaudWHzvg8keGwq14KNVhRLmYVB5foTwGzSeHChuungnc05YM+lEKsCq6kxiQq8wZeUgxnlT4a
zGojMwx1zAQ+7cC2Az3AOkTr+8Zn1Oxza6bZEgeoyDGjAiNyZB2RXqZrgkNn+SRsuBVHhjYZtOpt
MuwvtOgQ1WpOppaWAYezLY70I4OZUrffQ8Wp7e5lw4nKhl0cdDfg9Cy1LZIdxh6O3rNFRC88Kp1X
I5Am1gXRfoLOSKkk7Hg+4fucJX1veRBHXnx3XRZgV6v0JtHgrCK+DlBKaaQgIT8fnCnYtCGDOZyO
FggDot9lkCZIUMwcCM1/k8j1E8pYByHRlMUIwa5Y3hoBi6lC5FvCFggySZJSqJ5EvtlxrzZwz/Mz
2KDEOOy2dB8ekvdYhGughPyMKO6NFhA6KSerSQhIyXAL/nhFI84aidUv0LYiJUlrMcyPVnWNiRx0
5it/X3WLNlUVIO1wpZiyKeNWi6Gceef+IyjGSBN5UZ+0z9tYay329htOsMPuMLTRZFkRMihAfPwl
Fe4ZKYCWT93Z6GIIsL52WbnSfmXibvdI9on3EpOA3vnc4bIi/sSuEkUx6jkKxdX7Oyv09wl0U3Uy
mcFEMBUZ1nsiKGIlcvLyJrSJpaE2qAWrhHthf+YQ1zfku9uZWtt478Osw8IOUbrsCHbxJ9P/uRXF
a8sd/YWwFGhAzZHR1umgfgJomkzYVn/tk8jN0ua33djcstZ/g/LZGy3gsSSwqq+Z7pEsi2KWx4XK
K4zoo6JaXQL+3O6NBIpSmExFNnUg8kOrxWsEJLL2O5ImJnFprKIMe/7zo85t2cwfiesLNSoYQ6lu
r8ZFi1j+Iv+PVnVkf9lQlGL23foNCRv420qhgEqqV37+t3IWaT4cvUa0w2eXS5x0sPsPMPAPve1U
MDYWFlWmSBqJ52uDFLfA/jBll5aZM0F/CoPxhbU9Kxc9wZ8cxFgjWrF6SLrNTK1xGjrJ4TQYgFiN
8TKuC29NvBdKRsTS8eymIqpcLb8rNZXDeSALrktRTs5L6SPZQhNFT6HSNuaW7x1AAvtvzeZxwv5a
yCfLbHM+O4kmhFuWoiGDC4sPvUw8CkbMuO3tPR7RdN4Xw/aJy7cVOl6fvbGPKPgEmyZ63NIF2W7c
0W/sRVCUhD6BPqCQfs0WjCxA5BRXamglS6li5kT4CPUCaSCWxdRZg2qSMRtxQPDOjiFct+QDh9SI
auMZDp4ZV1ceoGORJl6wiGV0W/b7IocxLzr3sMyEKB2QsTxYDjT+6PE3eYYji7dM34ldDfAAQoD+
rOxPHN2Gr6xh8HJRltNijvEqnq3roqNk8xN0HrZ3+hDY+2x2TOxoUEL6Or2cgFU5BGSyDckiki/N
8CVHVwmpRIdzw/OU/yoWEwEdrEvUUgUEt4SnB92SYM4kmyo70RqZFWQ0rI0vU4hwAE++iBnz2TTI
gdXSJZ54xBvNxx8LywbBwygTh4ksgHE28WxQ4DXhKWJ4yWZpXv2LMM9GKZX+H6JhTu34IlmZt26z
YdP19aE56c33Bg7pTo82sv3bUJgIUz/4OiAJV6wwtzZnlBeyeAP7AJBb1IJV5jRKo6hKiJ5oFjf3
pevDDa8Ui26jSs3MKVpzkbeTxb2jxkiDpsd4mbf18Sw+KCnYuCZbznE5F4UrZg8GqYeWFkEeCJJ3
BWn9KcVyoidi7DZpFBAhJIsHb+ry4mD5NK5K+r/ZT+a6gb+MwGKbKru8c8PUvphDl/U39orqsuZP
ld6DABwoQg7t7i602Ay3XHOXcbO8mun1NxYi2vVXAy1GgRLML0R+a8ocJ7/EnFuWETzpS3vzMhgv
6r0TUxUQrg5NmGsKSmsM2PpJmsSc8a4dslPADZdiBIgmDrKVgQ2utSoyAdJO0cK6XW3oJ6Vy2J8y
YATqbM++1qXu/hQqA9ocgBWqbyBrVObJsSoQORNADwUjfNYQFBSwkaBfd/bglhh1QvdwZH3I1KbZ
Y7RQ8wI0DkRVZ1UizkfY5L1oUKE844gGVcmtb44xb6GJfMFklzewpgeLYYEgnnE5TtPnJGKwt+FM
hw83uNTx4KO7g7D8Gu5eH0veqxUI06x2a5gGJ0t5AGx60+45KmUoHVNg3JXbmS3NrL7fUUul2cGB
/7lgUKtOjpiVkNkr4Hgf9V1k5/xRYn6E8zhrOJJPeB5hk01+k1j3QvnKD7wf8f1kC7SArMzD0v4+
0BdmkpQ2WXxObVj67KBE3PW56XCmpxOY2kmVrXzvRfyAYdYriCj26O91f+0dJKYuJsgNyvKKzXy3
V3u4m+Zzn69f4QNW76HWgAerZLkU0toRjVjI5j8MUkApcsCFYGiH+P2Aa9GnXoS2KrARdYv9MNCZ
X2n3O5+bcyxnM7dH2AxBTKKB0/B2nwuKrwCda2a/o0HCLIn10U9Zuu5EtnDI4++5xLNipvX2iptt
Y+Yq9/cP07i8AwcnHxdz5sFufkEZxb98PC9Eg2M+i9OuRGWoKvBrVSdtkIWIBk3HFhfLMAw6B0Wh
hfBjlJ9QThyV1H+lJR2RSVYqR7I0pOVvIoU0CeIbP/wTyaPeBBbKDrvQ+xtPPkN7BSkWDNpU4Xlx
5NqSnrA96X7j2se5rXe1fZ5lZKCrmU3V8hEfoq4geKelyEr8jTYSr3RXaPGwNo6LROwmcWDFOOTy
zcuTnxCCcbkc9Aby38O/uwbI/90N0TQLo4KoHR5fqGo0xUEhJiD26sfi9hosb3Z/A56zbLiLZrNY
efYQH0+kujvo4ujWu5SJfDwghsv3IkeMGxuo9rnPivSHxeWo8HEGPA0xDPSTOGusoT2lOE3izAgS
Cu4MZZ1hLNRn3Qs0XKeuBVH4puecr1QZY3+JhQgQ09zblh3+6Runsln6zS1jgSd+FDTs+n867UqL
Sr1QolN5/lqRnaKR05MTu/dJqCzXZIU+Y5viJ8CYJagZwRt5bU7XSD2FD3gQ3DdX9Hloh/uVoaHa
GcSk45py13HJ3yoqCmGbgoOU3/L0mYhEVIjKALJ9ZqbdQde6TD4ipuXaLphVI0VZEnhyJ2tDrxte
LqsJ+G9hZturzeahDzSkdE+khqj/ukztu4p9WSbMwrDD4bq4zIkMrrhVzTsUMrBAXTD8Pg8gL3nU
X/I9y2wjWYCXOWnnFgTT3SQ01GH59Qz5xiSwa6Gy4XolzKGLpiD9h82r5n8tK/RtxS6yHkdKhowS
Qv1Yfh5bD7ygYIcg/eUnABvzJvAbh8LvydcAgc13kGD+G/PR9VLFle8s/VUyg1gih0mbduqMr40C
MFm2iA1Zgo7Z06ROPt7EKgHVvCfDufGKb+pyjVqr3tvVIUfEcO9jDi+9Hco/N02qRaiHw0mT5B1D
3V6Z62HjTGNII3/csBw53XNMY+EzuHnVsHIxYWvYLlcRp3n3BmBF65TSxZj6YuaAN5XG/DtYXPcT
G9DGqsHwxgl2U8kJd0z24fhjDEmZxkz7pgrdj0f8Z0W3EHhVmdgIfi6vw0frUSLY+HMSxXSYOU1c
eAtw7XHHjMBEjlD0/n3GPXxpjb9wlhlXuIMFc3jLhX+cfBhXxyeTUN/ufPuV4N9nrYpA1DXHsu1l
GvDxwFuy8Rxz9BRtHGd13Yqkig39U2fWQ+fNi4/lPDx0CDl3UD0AxI2B6l8xFxXD9YcW+OEH37y2
GvtDd8pww3Jq/zzQ0EoTaophknahT/QI/VRHwCa72gGo6zy8ragT2YiV/A0JlEfpDyzhprOuz/85
RA83Vd7EO+jL5BLKmesdddg9HwzIv6Ah1K4MOMoswfIb/O3QpMG7+OcmIxGOzhioIw8zeJ0UDf/4
YUT6phi01p99ZnTjZTRpmyxjhZykT/CPJ3qjgf8V4kP98iNFITzC47ZDHMrMO/BqncLXS2rd2sYT
bXIEiFqOEPuU7TpIdm4bdYJg7wVJMp5dIHGDFtmCZbVEgtwBvICJgMm4b3UReCT56Hs/puQfsFuY
7VM483TLklUFXv93PslHJZcBhvc3G6YnNesOrrVudjqNoANngUXBBtQ/oqWRm/xv72gQLiRPHgEv
hhZXmdgo8GAfPScBvJrweU5sZ+dyyF2FgyXAqibVQ4Wtu3Cpz0UCfyni0nXJi9o79zMgQTG2wbJJ
5JwCki3YBswziOPJCtIEfdENwZ1rja6uXon7g/sgXQS/YLQjYHPXgNCOd1wgtGgJyx2yKjZ9dRZ1
7CrAGed9uCgMnaWSWM9aehw3O4ArpgyKkQ/BAa4jZ1X41mV5prkTC60Up1215m6EJon3/on+7pxN
7BTyS4aRDbasnMYWHiVf5dTFl2xbnCgjHCmpUc0smmf2TRfhgS2zZRqndMkvHSyoVFczkO8b2kwC
mNw+TLOJWAhmhk2+JNGmmGCH799nXX6IDoEsSuPZ4zVD1uIuCtaI4LUBfJeI6DBW9M+xCRFbihkK
/Nfq6NHnRnVGfD0tROkCR8T8KLGrGoFdFeihFSJxynNWA+ok2F5B7PjQZXlIG39W811zZNv3060S
GbmOSCUdVPczgbcTcrabDF9td4BcEOxIoHHXF2w2spCjKvXQ0LxlC9YQ1PsiVyAWlix9/g+XZcYc
UXqXCWvxSyNma879CLpe0hPz9MITwMJiw+juhJrCnDyIL0enGATjK5HEJaxGIXIdmfLXmbCKhnMp
9rgO6r2EklfO4sgZ/jh6/H4Z/tQcbgZwh195p1OVIWNfRDamc8lKrbTabQQ41ZaPx5QZTwOny3bJ
ZwRI6XTzPI2du5OZ5ph53bHa8x3iAZPdtFjs//NtKFfSKxQyK6R4LZg3oJDYVgHVNakS5OGhlT3K
Pg9BEKn7hAT+JxP5AQllgrAshYmTLgnMk9W84JdQZFIGiSLJV4YsY1fQ6fYj1Mun+GZ2dPJfXizn
BIdWE38KJA84ZLF289qqTY/WmkNcoKUX8uTrHpc5MwDgp6c3221WFiXCxNveW2H18pL3ilzYSG4z
2vlbKLI6VvDwp6J0qbAbZyxXr6DIWyuMVRvoN97xeJOeh7ttPC/EBiIruygbinDWqgarV58owxAQ
HvNNZU/PCPftvCR/ZwOaxq8CkEPcOMIe5DYkIEL/nhf3aSXO1JKlieLxDPfiu0TkwAbrM7EUME6E
23rszW5aVJK8gqiwBLueJj0E7gRqokRG5rcw9nHfVmrAD8ZqbuaP1BkdcJVUnhy3pj9xmndTH5bU
TeaSFALwVa2hav8A2e2aRZHdGrxy02a84494AEztllegQMVsE/uBJ5menEWEKQKFXlpvSH0yMlI4
XDd+JcuBV2OQN1T9lPP5wLI7AK4dp9cwA7b/HtmHoyHOMZ5pqM5oO5pA+EMhperMw5TYPdZS1Kpt
PPwQ5yt96QV7QTF8/RZBSUdbkioIzMA1IUjV6pMGRuiyTWX4zoxmIG0v1Cz9EvjUQTEZaQZWJGoO
Uj1HmxW7ZScED9NjUBqDGRtSrgUkic2tIejdLp8i+lMpv50iFmoQ3sxFFHDComqvB0fVwJPl0FeD
sAyDnsnEd9y0UMAm+tw48BZA6ZvLfYuYa8OlOyY8ksGXaXRVXHaEMRqNrqkv2UDrZGqX0wHYXQt9
Jc0XxhRnII+Q19gtSVUZxuILtefwqV9oeai4Jx/1BPulkmj72HzG/YHuuPM0V4Op1/2hrO2SfKec
sdSLo4wnxKM2QaXm90Kplm2BoK+PJi1eFQV2hAVmNN6dsDP/LCQHNppZZTGf5DDERGaDF/gJuRZG
o0uoPhrTBdB/xB5P5nfTCiezVw2VatKVMR+qWYYT/5UgHlbzHR+ii3R14LGdidMqY9eQakcDTWby
MW53ZIG+++9HUXm4upc57+A0usOW7tAyFSOnZF3LR5x2MATD9I4v7ZCP8ZzuQVSUO9rWuKTxdEzy
wDpDdsi5KeGbhTodYot7aD1bFPz0Ubr7CAdwIuOBOfBsDTk58fIHI/hG5AbeLcZSyt4YudEeVtX8
1ZAbhIrGjQVeaIKQnWgSPiT4GmNMM19++iZ3AzPOsAPaorpwaOtiv2+H7Rxc6SYMoLGP6p3ItncB
TxaeqT3Sj54vt3S9culbbbAS9InzytGg5ZTHP6Aks6PIQSd2gSYi0pDdeJ4NwsepMg2ikr6wcKIv
fJamCbL6Ym/e2UhNE25pkmCANYfqTL17qzQaTjwiKfzWF/7fBSXKv1hdj78dgbQ+Ah+P8NJeScPZ
nq4OYKp0b5AcOUgSw1fimEI1VakY8bR8ffLLmxaZtUCp3SwuD2SoPNrD5bg4UwtDU7wh1w+MD7iB
hR3eOXhGFQ9JiiVrP5V5ZtogfY2MHW+9G7VD9VKXLks2Xko+l1Ciw1W1vfc4g+xNMK0ahL97T5ef
lW8ULsfMVi0Y12XSt0QgX8s8BbTySxmun6VV9ifnyoKQIv2vQZzStmHqGPCZXeUxTkbB0FM9b1Yp
EWeOCgvOVkeeiEyFjw5uPLD1O4u1eRbPYSKzmEmoquMy0uqfZBq8UYoyrEJdidYeQshMXGaMDprH
BbaIUf1Djh33NzelyNC1FfgRwerhu62EpSF3AZUkZeAWyXBVxiqfnzLuFPrUTkGeo1noOJfhkroN
JH8eCi+TThkjkuw/Fv/hdsNluAn3gF8I5U6E3l9s8W11j9JjzkIUKLaCzPpzkgkFucaLYySNRXN/
S4UhmZEtZLQ9YLaGKk6/pDV53iNYHBfIs5F66aSoe7qMpE2VHLiuejOkYncyNXJNRBARsDVxBbsX
U2RWUwV8VkzB8cyFPzycaKhD4CY+KE2Icq2HvrMd/f9UGx/5fcldUDUNKS4G4njdyvJcdid6hoeC
uqzecTuaVrv/u2YwmWCFKh9ZZ6B6+1OibGiq5ZtCaLRNr/XBVfQCxh4ATgrrKbuVYoEOYO2poaMB
OipYhyDhPlw+63dqA7TalckotFR5NnMOmgm5YWKUmuKtzKzJRzNlEffvsBha0iOXcAfIeBxAL1n/
YoRfCpL48C/29aedRu4FT9hED6UVAzpcK3RYKh3ZQU0mGsHUJc873pqbvi4Br/H+coKIc5EYyIG8
czoiOM6yp6IAY8eVt9nuoYoaIlJauen+vntNUNMdKebAY8Xn5xuUEzYz23uQk0JPJqpnPJcvo2/e
MYpQxXORRbAHbw1QxllgzxwbSwym5LjKYPKzmpLpg1NhiX/3DZUHq7Ypiy3lGNrMUnMDiifOLUK5
Tsi2tl4GD1+7+xvnANm+xnPLdmpmK5WDDkRQnImTim2hr1doRCXAW0fv3Q61Qraw4tOHaofzViQB
3z81pR+RJnIYloMUIsIiT1KliJtT+607MJKDqu30xBmKfx4pyMIAt/VxCelB20n6zzi7W6YWJLCx
GRtv/fabMp7yMyn9vvY/cbSGyxYRxT1wZskon07dma0Q/aYdkNltOfzEwAlD0oXy8gGtfEeRTRG8
qwHucoy60fGmmBfcNj+/KltbUgKIDp7JBPJNq1J1+6vMlSSQLD4E3lAkaS9W5N+Tomyabn4Yw7g9
Z93ijR9/UomTJ1guRaMwMohocXP/F3d5WfMvLtg0Dva+UzmWze3B218PrxRWYFItEzCQZEdkzauu
+Wt+o/1G+5NK7xRu1oVETIcuoZUT6NWW3DHDXjGbsIk2R6RqsWmJ2eqkoghbRNr8Kr5jz3vNYBfC
G55C4OoDX/GNd9Fz9qn6KLpzu/fIq/Eo6/urfkOoeWASODZ3CY9RNBVeaKtlOQavK6dMnEejjjKo
9G0uHcgkvpEM5XtUnqHTRBXUzZme/REnjp3ZQKJPHr2ZkrZTcQ2Z2dNLpvJIHa0008B2UUyS0N8d
nV0BnljKd/ojcDDGvdGLMJkMoldQLzqC/1XubPgRPQzKAUo7lOntJ/i043NvvzK/Cin+2s6uPkcA
EOtIUk13lhHrVSqQjl8ijk43XQMZY/lc2y1c2FaHrl5ePvRhD92P5KWrW/L7iFBxWn/bnzendjpb
JTnBXAMR5eShG5OOoos216q31482lcJPbG2E53GmeFV4dIN3mJOK7fArU4ixIj3ivedLUtJa3aTj
uBJD4y7iVB7deuT8D7TP/NYxSQrsoMaJxQYp2KQYtjzBSbRyOfvKFQdjzvPk6qr7JRuAnQPHj9lV
ZqvTGAQhTfdUGJIuerlHgKJ9ok6LpBndEnN+Mg8hH85FTE6HJJlxRbjJNUv3mxwCy3QpNmCLQpjH
uzyLQ9CiGhrsdTiuuvGpFJzrNd3epMl1m7jjncsjK7RC9EeqYG1A5rkz5ZSM3cbTQ9kD2VDduW1a
1slt1XXE40NMD3m4c+Ajiby5bYZObzLLP36R4msAHgZPP1O6qH0b9ntjTa2yygeMiXls9IDwjvh7
vldfcP7RFOhmFq3aC9hIrA5rpoWrN7KeQO61QmVvjCiBd/vBEHAUXYb+D58k4virotjAdB/BMsMY
/f5qiTChJWq/Le0oVVmEy8rlxUuJz+2eM/YPEiy2+EqqG1YClpXTsqV+BlOnlpPdwsoZS4a4oNaX
1QoJoGFuLbb8i28AcSX8r6+7MlqfJ4ehIA/E9VBTTUNjY8NGzfiXADkY/CSo+0Du9oc8re8uNnmi
3ktWmF0NhOe9H+nHJIPWv/5c0VYGxYX0R/QvjJ6GpzCu0/Y0qGqbSw7VJR9vt5KinxF4cpBrD5a1
iKd67/roig7VK2/IcDvL4hSe7vdk2ANdjxHLh390V+evIr6jQAtddpG1QbUGYVfJ6dzzFuZ1A8QS
kLMVoUIt6bVHiqg2UUh6iomQw+3J2bupOu/B627JFR6dSEFnyrZVlnE/GRjKM/4KSld2ORuU31AC
LEuFjUW/CchmaI0nHnzGv33EerPwichxpzXyJN3ZtA6PTQa+sZa14K3xZC7X+kZ5ImXIJYN0GKAZ
OiIO+s9hymSJM6PA9Y8hedLO/j/5fnPesSFSjR1/6UvJloD8xQcgquoH3GpMxRimWYWFFNNwTSD4
DaPQ////B9XJMABdQF2PEPRtQATi4POE8T+3vCypNWYwBtUaUKpOLoQdtJZMieZjh+cfu0e5zQyy
G90Ewgm+XF0dBg1WrrErY+8X7WMIuIoSvlsLAT4BRTCYxzOmDNazij2NIbJp3DC6fXgu2wQxJpfP
uXv8SiVIXZscbmHaSsYTqHLdznHoXx4Wgy8dKe2CCXrdHYMFcozRrfriSr3+6sCXr3t5CkhZ2Db6
aXpbLQ3pIFX/OQ0TG9i5Cy3PI/w5MAWSHCckqCsqrzMTdSgkUt28+rTsVOqLkQvomnYaYsZh7Glo
L0SeizKzjGeXNpPbscbj5JH/YaWh8nDES3f3coBEeZHEcABx+e1H+xESuOg3zb4YFz4lXfLBjXaD
vnuYLLp3glFIK0rZ3AY74lUw+DCNC0iS8hy/UM0VP+U5sSaQ46RCioTNGt32uL9eZ5BwaCQ0hreb
XM85uom3XQFsiLSIetd8TyNE51wjpt470lPQ7nPnZCaeo72HP1zo1fqs5ce2Ox9EusS/1INxwKSe
GwjJllkoB0EJXsosJVfJPf4A4VmJTdP/yzVvZf7mY+3zjnjLzPs023s/vSvSedH0oly/mqb0q+hm
f1HVGL2KhZe6nemVN8NIFFjwEQcvBMQf+zmPldjnG8GCLwabYyETAyiOndn8ln/DFydZRP49UO0Z
8MQ3YZn+y7p33EZIdm5rf1aFsQ0fK77P3WSGpvrWM/9x9kqusS2xLgHrRuAg51Wr0znM+siFNM7L
79YUFpX2S0cBiyoyscOkAHefPSw9KnmD8s+nL8JzNWxi1neDtIDTRJgNIEx2w0cPd/tldyNCBPQS
ospoR8FwCMbPPXQUYkvp6bNFj4YiiHuF90TXrZ6GXH2U7RKNryf/UbvXO+sBOUir8GCKhdXAR4oY
cXtxn83qGRe2jIpSwYTUIpoi3jpyUFZ1QwaZp0qg6h8sB3/bJDGGe1Sm1wqdMiTYN4YmACcsJIz8
I9Aq/X+wQ2UG8kyaDEDMpd9TBwm9737bVbCysuLnGHx/wnBah6gyu9pBL60ukvZ/7upT72G3MCtU
D/Gd3BbmSny0zs3ip8C86atAU3YYwVzfzxSo7Z/e94Cx7pLgqlfJaJZNR4cOHMordnhPhSicPUYk
+EPKT9lQZoLUncs6qiu+MBIUDuIhs5Qtffk5pOjfiIXHsAydSx3yhTFNfFUwG2kQfXxhGX8c4A8N
CJmFXZzRghqZaNf8muSjF166zhMdHZ6ZY2DF9ZZQngr7aSw2Y8bUe4tmJJP1ofRrccJvYQ0TFQFG
21yN4dr1V9vAOKSskxiZJG+os6QePhDiGmnCAlDdPgAqr+Q1k3X/rRxL3r5kB0Q97zL5wPQPg93y
sbpo15rRqFyMTgnoUlNFz2C/J4xrvQbB57xGtgiVQ7ypOrWRjWfqiOyPRt5JvUGSQjhSZ9ZTPz9c
0Lj+Nh2trdPuoIZUu69kDG2DcKtbdnAqsIXrrL8XIvSky40m3d42dnD9V35FkToZ3cu+e8nA/4TW
C78BEQi7WXuRbj4ojkt88WBrGBTaZJ5bUR5AUWOHpXbof9uwLnMEG4pBtSY/p+9wMGeq3VLvEGQ8
EyeNvBuNvGLYHcJE1Ovkx5MjimmlAg5671XL6BT6/W4TnP4yzFigtqu6bDnp0dVLU4Ph3U7XFsOJ
PVaR5R3Y1WlxVNtXwbyV2MeW8mxZOlf2biamPnmmgO8Q7WcFew8IR2IvyF+fs2UOUrC2n8EHmzj/
UJ+z74CSENI1fN/LSALOXrZn6ZKZrRy3J6rUIfwzmYPp6tz1HMNzyy9qjDQvYL9uEokipo3Ra63S
fNEksKayjr6WeEtBTFDsoXh0/KX8qlgDguaiVWY97ITcvjEAH3gaMfP0K3C6Df+iJx+uK7aaSQSQ
BjFyHRmunOmlVDD+axpQRwJdj9KQmtiLrPqXLv4EcgGDue4DJa/Vr/k57QF9UwyFSuUJTUu4MRmV
M7sXrBYAgRSLlBN4EWPcrHmGXDJAiC0GytvYx2GpaftldyopVzIrcGySnP3mL/V1lRfyzZIi57tA
Ez5dyAb8/XI+ANZLbY33fbn6bgqbeUktRDDoIkDjVjusUix4xbnK29m3pf5wVbN5OnP+Oa6+F9Kq
OUOQXJcjS+t4a6rtO8SXnP1kcA2xFX6bfEHhsmm7+Btse/H/KsjLru3Ozc72CuG/sQARjRWgMqQK
rEBMYfJXAhoqWaErKuR1AqRLwh3PjuzGPjAFBI5bAtnhJa6u+vTAg8FzK4Z1L0vpN2YfgvOfhkyy
bheKRGpmLg9b5jN6lx66TGeZuO+eSVHqhYCw5hj14CE10LqpnGNOB8u6ALNBaQ81izXQQzo7D2vW
1mF5BaHlaAqbLOvVzalwAoN3CIkRuoXAzwrEW0M8lEw2xOuDYAp+G/yX385uVQFvwUMWValPMYiJ
Dc8k0H4hF1OTnEXjmbU9puR7UNSKCYqfLP5FVINYMQkELwSusgPPOe2y9dIH+gu5pP6w4MkMEIAs
Em9L48DVaZjbWti2zALCrRXyx5fhP8gz0Bkte2xpCsAJN4dKo6BKws72U5gir+6sUdRG0JVgE0w6
KziRjlf+5r0yG2DvNFykA3WGA1l7eRN8xjU//weG431Rtq1w4RfvAtw+KC0kmkc0V3q+ktiT93/E
litHyUzu2EgC0afReWtcX3Ct4ZNw7pxRPYYFs2+PAlpHerTVph9qtewdfArKzVci2hymdCuj+39p
Hk4fefvQSeNoueiBomDa99loFkSq7e+7+JUJhLI3zuYsXbGIRWZKZNjWC10RGfoNMunTrTH0elne
sLzBT+tyewb+xxlucDHLMAAO3AxKlpFoibKZToT6KhSKpTIEtc3zqHwyP8WGHHg9hahYJ/UkOAXM
OWj9cpSdLawHSRQkEAPuDtfdSKk5wAUoseybqJs+HbsR9NCJDGTSNU3oBvXyToSEaDR/PhEHGMO8
lePXKqjhm953hmcnas/8+AxZ8vq9f+pGofMbYHF+kRBbUMRfdqpwzFO+ir9C0LNQ7XLjT0Fdxaqf
GAKONuioJrT8V7oUBodzgMOLN9lk/pI5zpXUxGIdn+PlZvB6dOSIZFet//urhB119vDILWZzriWR
iQdmib0CcFbO8oqOdNOTW8zZLRwYdnmjscTf9yVAAD8RCy9TjAsmQKKfr95JD6cVM+CHsaQY2Cem
l2CN2xyzNx+Q4vRDA3o1cbtHWp7by/xngxXpBsnvvNJUabbcFID+XbBTdObWMkYhdHRAiZla/A7S
z3CVrcmL/WPREXfwJ4K75e9g9mGYjbSkPwk6bwdy5eWwimDYmQjfWSWeVqs3bO8FHEoFufXTlUme
1G3FkP8snfyaTsezv7TAxFRPStigNzVmeLS/LrgC2bSG1eVIUnbPekfK1DAnuD3KeuTP/ZhB5LE+
ak/LIGrIGOehjy2jDOMbUL6K8Q8t1TyZqhILnGJbPutA22JwDSsIIT+yFhlkMpTvrTo/AjS3A0PW
mG4NMw74Qd6YW7jjSRJV0XR1EAh8IOGmXIBbHva5NOViqXQqX5xWvwYkEI1j0zls4BGk6pKE4XVT
RUUnTXOQYq8f1yqTFrDrGJL6Zs/NTCV+xkZKQW4z0cXlNfBx673+vYLhID9K/PBPStKuu5jRVSJc
fPcJwkq4YxdwkCEKIaTNQ+lvILzSCxCeeWNTJPovZAZS/SFxb/DpS4hnJX5f38fiZpDdibSwvGXr
wj1qOQ0URkIrL+8eUEwgUTEe5gtsCYzzqrCsxRs/6YZIZu4kaFl/e8vUA+SsviuS6oHOUTPKnrCK
hwwLAxEb5/qzxdNEZol1caIXSMBv78U6jDuAr38v1f+moxO3r5Y4T8PUfCqO9TTJdum8igrzoF3A
MrdEHiBZOqJtycO4aR636qxj4hoqdgx7kVKXu6DCJgWZRzwIuRTmOKgKqDBMOHu3MA+/gJZYUbil
BedVbrGPksdcvJkcHI9iLBwUJkOMEknleTvRPUEMpSIn/bFgbWTOFSBZq2xQ0fpo5KLa8iHI8BrB
Fpdzg+jH6XQau4O+C+bqFAsIjWw824DgxrhF2qNFsvq2e8DvkK+Wg9jj+ckVmsPilqKKRfmF0QNU
+9PvDqypdrejWBxfzHy6c1NaEcBguLGvEaVmQLvtcjnFO5YmVPcW/OEwLTp3LXb3TcEGkmefcRQF
+9FmKuiF7R54nuJynPBJ5bF34n50ybi4YjHGwy0tLTxRMCij55QOqKqbjwLRMt1JP7dpyqmFmtoq
L1hpq8z40DQ3hxnmuSgcuDEv9jU0iUxchUCZMkP+O1xzxinQ9aOQdDWqrSYdOudaB33EqgJgpHWj
bb9OSvMTF5Cn3rHjKnGH0T8F4rOUaS+/1SqG7Ue/XKoNUE2vxTU0K3Bknn+7RkZzmbWZT9JIj9fp
PRgqfbGE6iMc+eyJYCLX1XV9F6Bm1F5aGeghJHzKUVJBCVCYjyXR8Bfg/n0uS+sQHhjtDsiWh/jc
HGs5Ov/gPCGGfOBMtVyksMTzn6XBANjr6oS/JRe/PvF+Xkp76Pw40b42NEs9JxbjNvfDULNbvHQj
lJRAl4HqMjn7P2I4F187SdQah8LHPkEpHPIyYC7dRr33BcfsIAfhGUwNKQ+lyDnvfUrtMB3nTloh
8SKM7mhMt3qT1qNTc9XjopQxlvyCdYbNCFdHUpG26PMhMwVK9XXpAYb0E1d8GmouP0NFDgvI+8Tb
SrgRmvnqWQjqpJ0rVhtaQhg+Z2sC8TWYRVgP7MCoaI5UW9iyvHFXCVcFUnmS1WFECWw+gabx1GAe
Wb+aAniQz7y+frLq5fbsiT0hwBQ8VX3uG6KOuZJXAByAqFRhwJxWfdBl+9PR57cqXvWaEeLsTbhq
enomPDlIvsZfqzCsbpupCE68utYDIIq38UOMLAm3Yc9iatCmn0xi7hINiEIOlUaCjdmoAWtHpu5K
G2DvNeHLu2bIHTHu6bXfFnzfZ8y/Z6Jo6zwCi1jC8IqPRXYWaXyOY6ZAtteCH2HQ1RHG9IwJ0ImD
qkctlXJGXaq18OZRF2iYV9oHACCe/Z7HezneVjhQ1FmNJp77xA0BAEOzaD05SjqGz2f3fZDCJ/KN
gSwv+hkFgf01sLSTLHwQXH3vZl20RWmgTZyXBPG0ratukBe5xorw4KTIL3HhnZv8MT1yTiw2QPGf
r4t3TpxMRqY80tpQDY5LlAYTg4H76sSutn17v7jAzqwAbDcrooUpLtH4hshrSeToUfiwitO5nvBU
WntChr5gQfL8YqcugGyjq7fPqjYa5JWnGNl56JsFcFQdFEWsdSe8japMPoplMik/F7C30Oo0Yf0l
TKcuwuuR2+DuHwTYswTk7W6KQUdPgSI1S971L01Wyo2VA3NRzIUyLXr4/7ThOzVtv5M2ZSydp+gI
C/ffaHDoY+dZutY4/gYsw1ggccIj+i82rFUittKOrVDCzzU/l66Ah2qOeciYXl/P89+fjaGVGvXr
htLW5zjajDI31iHdTe342RPWQpW+4L6CWuMXfYCZ8zIJaiFrYrx+I7quW8d3sk0zj2AiLPYEKSj3
P9sNNa5KsjMimueWSmDDphExg2K+ue0M8f2bFRi/RWXTHopHYMXW2K+hS9LwDrQ/qPD65dG3JQ/p
omcnlYlAO07N41VQWv7TS6ya8NQnfwSZzg61j/QMnBrEc0SXicPOrwMwH9fcmTAHttR7TMQHzAIK
Qh19A3xGxKr5xbhy/1xBmYFtWH/61i6IUhAqhVDZQg2KD6ayIC/si9YRqbpW9yvy3gzqgI0jpNUz
t9V75Px5sp8vPvCap7sYXm9EiTwPyGfhnKDhItv1yVUZwxTEYh0vxBzF6DsUrI3cupDFYKOpQvFq
DUxI9VtPZssxMbPdkA60MDCK4wT9LGgAm6CSNqE+bET7So7Gubs/ZMljrI+ekz08H4hVNuwqUZjM
CCEpuyh/TikWu23vzHm4zCyjsWhDkiS9zwuZQRnvtZdiVxUJ2tyR9M1Uve6zlvY6H+j96INXsFhR
zncGPoQP5ToocSZV84fpkIvLd1cQcw9aZ0XkkPQYj10imCejjZ7aBcbt4lAOCKeh4v6wsIwyTW8S
Zb4NF18e7cYHvZL4lmGWyrUVDinArXqYHJmgRVOvHQw7cFXgH7UktY+BkVl76W4GT1FOgL9HjkkS
zUWgOXG8NOKIW7Ht7njnF5Vvq04Pj7ZxfWZ2GlUrS68yOQ0vB6Peom1iKSrE9aWtaRuw/4e6c+EH
wMzjbpY3XgLc2gFxt56pCb7hQZeKQetQpVD9pOIEQshpcJbH3Fl6llpDxjD/HFCXeWB0pE8QtKMB
ugRghvtdkv7ZFf2sI+jDPMNpGp/mG3V9SDpf7bXAWLyQlsDxx46Kz/3zPhMOoPcT9Yb7BMzFbqma
NCursA1s6Rlax7fuqXnCF2VIamDQhPKzR27a6HUyIjEzigvTNbsodYDfTRhGkfGACg/hJxJZL6iu
yaRSoy0yjRO8SAfgfcVhqEHbdGrzUksjW69pROUgqUsQlrdoXFj/ZD4IVvkXrjIguHwK1SWe/ygz
R3C3S63H9sHmjEfwPDAwKSvhf49iU07zfjOSvqJPweAGUiWTgyJlWXvr8NXop2CmXbQDqLhbKRjF
2Tt/1FDbzbcgCJYoo81HJpG53WsADqUu260y4emnpTkR7mxWclUd5rc9zEyRP6roLrd4xO7SuuTA
rVEIgFAvcJ10aj5WYpcFGDSv8xw+1iwSwxnmD/anyW6DZ3mA+kwMjCqAzyZS3kX3FknMUVyaT6F4
v013mfTIKM8PHcYRXLiR40rIO8oI9YgZsGxxCTQWdOTNI5hBD6VK9+rxs3L1joCmfNzBabCigP/e
yHj31e5SpFv5mR5hUoAIH3G+9QPp006x4xzDAIHFH6JYezyccdzYeV3LxgG4F7QZDrkUgKhKvLj2
bzYlSx9ePNliF82f66GE+la4yebfMOEQ7c8anN1vgFXE2gsBCRTSZN8s+eTjkJYtFqEM9hc7Yw45
m6ZjCWMQ5FGP3PCpSgyiEOXuKuaYc0cV5yTfujrpW8Ji5n83cfXD8nMyMzWlv1pphHlUNAhvFwEQ
aoDH01Wxpd9nm1GNNJ/7owmDDnjVlv5a1vjF/XRkHJNicMZ/3dmmLLQR31Y60Ix5F04y1iicfPRI
oft1f9ISRFT7AQd72sHI9vzSL3/5oflaA5yfaNrtR+89pewSxZNaHr3RKkfni7HZhftXV4pf/LGt
41Fzb0Jf/Isux7QIemOmIzb3CRcaxj+iKHk5kwd9XUCFQbcQlnNOJ2GQgwJPWynZiPEwB3pFNh50
RYREzYKIt7w/y+/0Pz/c2jj4zLBQ2xhDhhcFg5WWMDeSwsdy/z1MOjxu4Cqiq4zSOkAQ9ilj9eZZ
exiwveylguM7wMpRzUWNXqARcZ0WSntyiEMVkh7EwHdV/VMdFYpA7LJt5PZ3UfOYi1W2BuKdZgzA
HnvsDp7UUuBCehF0yn8WpHBM/40XjQd1T9ltgLLbUrCvujhl5hb+UzIWD0Ms9PGc3bv9aLQBqHk+
7rCsNd+VmSHnTHsTKLuXxARqMcGlCTYtfqsENWCM/5eWL3l1pgww1twRZ3GWIbKffDAEvEO8jyNL
qmYeg6P1v2UNvR3C7bnhTJG72SkK1V7j/neSh/RLVI5abeuVo7k2b6kSq4RQ+Mfas5dD3sB1sktF
Eoi9SjknbsAK7HwGhUjQN/h12S21Iih5LRoR7IxGeF+mlG8wjNCVk4WQtSmNqiznFexUEj9hUnp0
g5JhhfeeoSXjAKR0/xA3QQ9U7XOcXczj4frjfQwrNKYwmLOeqHWFFoCI+1FOfq1Qbies38tSHzgO
PifYACRzLzgzb06n8FPlY+ZU+Fk2PxR7SHGyqg4NfxqcQXhdhaye0VZVaurgOG6Clm83H+gpeJzt
vM/Sfwsfzg/S2jLyZFRAvdNdEVlgUwYRbqgpTGR0GwGItfQjbMAV09Fl2O4tbx8dFOEqqlnYpQgF
IjP0lllNfj2ZmCgSzrU5Xd1gkCaUdqzvwgR4GHlXrRpjUIOw7dzhqNIbvqaWSS8gers1zjpprvOt
BL8wkPIlcEiclGZ4pwMzDgptB+n5PjgKfBphLZWE55Qx1DA1CBULGqZhHSn+KjeLudrNDttW2dys
W87632komosb+Mt2fjRAmhCPvwH60I8QYdc/0z/asjop25+MhLVPxiGTPI/Rii+F1aObp7/OeqPt
rIyjuJjuB1NGmwPJRhIXghpI0uoXFl+cN2NSBWQbJIONKv/A4be5mMVC1vSRgcqgMcSSSRjSBRul
srRHvRSTSiQ1won6iWakMI4eBKx3ZcyAfY9glmgyGae17BMNSxF0X8h/UIHvDlGWzmJHjCPlX08S
rEJ6yujGYIqph/A2XBso+/sX8L153pIAj+XJDARYqqgjKYd7eNu10TB0k7SALpQXdkQBSAfMZzDp
qtstYQTemDNJHWozLnYMf4Tr/FDlReb7fG+x20ZDOb8S2EGtCF7MO8eKf6B38YCcw5D08rldQDb0
6KMr3Xt1WfAvQrHwl9m713XVZRmKcJPHV4TbJW9v5zpPyU4AEAxr2fhsyk1xOKjs8LFcOPfBAJc+
peg1zi3Nc1UdIAMQwSMKFJTjWYf3pnTdqWx/4M0uHrqIvAM/+8pvggsh+325aTrbXJQc04Ga6Hsh
AoKhB3QO2tCNpD0QHa2DXKRJk0Z3CNoJ5yQ4jnKV9fu6pLPSmMoLJO/Fow/9qX6hwOrWe1ReG+w4
paDM6RRMOtxf2XBgEipIgn8Z+oYDcLbbRiNdIi8g2iOy1Y1SOWxkg0QrdIGET7wy6LzJPSDGKBJL
/OswsBgdIw3+bDXOOgWrbEI10QjST6jbx4vZhqLBSnat4yTwnkKk2XvUt0EpXuZwLL4uTHVXOfVx
j/p4q0pu7Mp8dngb+25mWoFqno/7a1+uhj+x2FHYKBqMaD/7KBmYD3JLU5BtEa5e9wcLS3TsE0oc
ld7jOE7YUp9YC/6swswm9IFSr8cpltyE+XR4MtFC6csazhAJY3FmM6r6Ci2SXg+ZQ6DyQx3FRtKP
gC3Rn6aazBMOOBKHm8j/O0HEB6QKxvLsQ8FWp1yKvOXuUcPzVD1jYGOdxxLSuSS3hYcXEIiYUuGs
MatDilOQ7PN+15yKxqR2WG1J08C80TIVtuTdflu1cp2vJDnnyHxdxeK5W7wk+8XIdrq5gNcKcozm
1hkVruhDt2o/yxC/FVoW0DtYnq1D6jHfih1jVwwhknRhfNDz7AvP2lF6ccsA0aAToyVlzre9rXuN
3siznsrSjShRrEPbx5jGtNI1/im7r4PU4ZJ7qUT7jQl4+J/C3A11BZa6VBPuuUovUVh+A1GmZtP4
oxTTjyHhInUfTMI4P1q+OleAqy0PcX0rarXDx31V6oWJU4uwqgvI0urJvtcmalgR6gb2iI/9WbyG
SEs890Iu0sVgAofrQHUsCcanaRHlhEAZZhvcFfuftHp+FxaU295i8RMNw4UKC1VrJxM/NZMLk8EO
Z78ySiEY7X/hk7728GzKWcERrkRZk4Xq4j0CxsCL2gdQyMPETIqhHPVZG8fF9lJnjZ29can5oLro
IOw08x7y9JF94tnwsoiGlZHZkmtINMuweOIvu4WR0zUzqBSVCcxSKH0xJykoYUL2wrc1Fp6ZbR7I
qX4fThz8GEh/dx/Po966pr21z7OPL23EtyNcJtspf5y/YcpCJuJAGLjNmUSaHms/HZ0T1Yn1JyT/
H1+BVk1uCzbF/27YqtO9iDhXOLRKIqMigeYuhxaFaMAAp+lClk9ItxyWzSZEmCHtqiucWT5/DupI
JYAs4gc8SJgdx/IjAo0elzhKkiooIIqjsBXCvMqS7IMjTou1edV99Zrfr+38vSYQlKHljpOS8RHV
SlorExJfOxk1+SUH4y4rjrC4y+n3OrPaU0OyXbr1FRMrtDNBNpvWNq4lPw1czA/3kNLqcCt3R/i0
nKtM9QisO22KWS2a8CRhqf0qsK5JTfmH9ZBR4DZlGbxaWeSsQj+nPXIRE7oVN/9gUWn9tjXQj9z6
yOurs6rS9ThWxd2g3c8VxhUwevTcnkieO+LYloCOXuidrtSXUPfx5gqIjTO1vfy20emHwxAb1gPd
gstaGJ+GVnNaPUQRGaXT7UDhq2BWQwKAXNfTRyJ91E2iu9I/Pc6hLtMyo26PeTOdSnY9nq3nF3Tq
oI4HJWXK1ODEzH37DrUdm3ju4wVj5w9jXw4N986g1bP6Xt3kUGQth0V8t6kloj9Eqa4vF1KY9bsC
uaY5kpIoNbnwlf2N7A8MNnYifiMmMFXFhoN7bTpirLIWQGIbhf7LFfT4vG995vJUJVUoyn30yix9
WRRB4bU2BHPjpE0/aSccQyZt+Nff+dCplOdYkWdSV/jZoax6D2PYEXSXLAz9bwrZHsxKXfJ6xnVp
7zNRBq0irQ9KzVQVfoLYyNyDQBXSRJVh5TpbI+/n0vWKn2ETdAUTk+brVFnFrHkDZDQDD9VLum50
SPadTGeSw8bOdygLgf5FbJQTI1aaUNNDNffkrjywlKbedPyFTOkkd5cLpR8+trIfSjWr3cWDUnJy
XSkhWMmTFdaHU/Z6m4ArSS+5CDEYoRC9AznbowrlEEyc3HowdqnV27HoShU1knPwPzrA8B1f7NMt
6LmMq2YuAziJd6gzEIE0UOPqTBmUDVlbYmSTSlIXKmUAgVJ6nROSwpyW0azVTNV4EJhlIRfPVr5u
rf73X0vJHq0+vqK5Q/WCYJeVE35/KoMgYf+pxIdqIyEmWdj7NUQcKlIK9u6QVlYP8NYmMDh3GaPm
nc8e5Eoiy5KZby3R7xcl/N5AICKpczH0QGhRc7jxUnPmGObDBWNn5UTZCDKIhbe7ITVIQ38FYO/h
IM/d84wi2H2cHAKjhiyTZ17zA5R4VxQSwsAqo1/YNL/mwqib21dMj8DgaqfpjoxcUUhJpmRAhhVZ
ApHr1kl2u6JHrajnDbRAT+J3Vgl5wIQh66Y/mbSPKIFEhNH+I9pj8SZVvHxqUVeQVMm0xVZbDiuN
q2B8fWkdHYBtDlxGi++Pelh3xFr9/EX78It1JOt3qFa854D31BuLJlWaHkAa3lizVIrCy9D6LeJx
8lka+3spHfm0AmZjJVLp38++jICoUG0NuK/TdTU80kvZT+Q6ph4AspYHLK5oMuYO/u2JWjgBDnML
AjBMNjLiFO79aGfnenLuZdIxTS4hUDDOAjKGPa1JBjnvZlWKE3IKz2Dmcs7cGy9LaVgKuNh4yTqE
AycDsT7OxgKkvFPOPmzUDWKrH/2/o7rYt7JEG3SOmpFmKiWBVZp71d3s0CyCj6iNy/PsfkyeWQzQ
rXHPJasi1r4bcINrebzEH+njrXNmTB/QqhZCmhsFsZbIu3Srmr23VfsZkkzDUCdMhAysO7S2FIS3
SrCJ7UsJBVpnDTjg086nzbcYSSXkOVv1a81yG5qY094zMGr7ssqfXdy3ZU426gmdj9LgUY+KdwLQ
/Z2Dw/erE2dM70WHx7LSmMsOr7yMFOp/D6eBGCQdz5f6z2pXaWFuUp4okzPPrJ//khK9UlmBetnX
WYXe/XzocJ2DfbkqJG4YA2dbhcoaCt4T5OmA86At7+c1IvgFh8Z5bLwlXVw7zTsl6BgDpog1qQZZ
OnVEsdsZOiFusTP+lvzwJ07+/WB8oAFxStPKfjRs2aTUzW65FX33ms9oT4ezaezJqbnJs2IO2kXJ
ISgFyq5DNhuXZDA1IcIioR0zE6G6uhFrREa89s0LM/AKrYmPRa70Cz+98EitTQmk6tCGXLqY9gKA
uSfyJ1nW+AmeLmlaFViEGGiIplhBxQYZ7WHmX0DlI5SWq99sYTL4TepxmU0PVVFwA9P+GqU7DJsP
DTzvf8lEHLKTUco4THKz/8QM6mX9E0mRHCpS/QImxpgOMjTuthDzIBW2tG3CcB2qcxpHAH0kNPpO
WncJvtI2Htp7IcuWGLmtRKSuBw8nEEaiO2s0gb0z1RmGqO2PJnC8nZ15TcYtvhnf7vidbg3vy3lm
bthnRaImqUKXocdgP8gPH9L1peUgFgPembk+hy0ku8prie/Puvmy5uwVE8H7aq/NAnfAoKpSvKTj
ttNZQQ9dYkCmEDZaNGDDr+IzzyP3vr+NpDxhRwbE8vY9HLQR9Vrh1N4YxwMRFh0Ba2DHRjn9rvXg
KoUk/LM0iayG5xNVmNgOC+NPzApQMB2q+2QRtoJGZm45ZFiuKc6rYhLt5lVsGi7fNz9cbgSMMpQ1
EsHiTDRKIE76oYvz9e3eL27E8kDYF/Pu9UrwU+N41wPopgYqIIwOrEnfaq1kUoWyXzryNNAxZjaD
h25u85hJXPGg11trVzlckHC0LTEmheVYu3Nd2lwTipzU0DqDUZ9V4IDDhk2MuiDLNf5BAN2GZyg2
avxOPqcaMCoU3Ei/lDC9LwW2JwXWoA/pK6lrJ6JD8lDMqlf+Zp49mTP/5rGYPRBC1CRq3VKFE9dC
t0AC6eAstV166jFs/C8f8ulXDoTNRckVRqYL0Ub/z9nJKpEXxlTGURL6AfAdjXI1cGXjS7ICOPYC
fjHGy7MfhM1L2rm8Vsnolkv2lzd2i/WwygnFJyN5se9EReCwRi5VY1/EDLTaEhieSGYaR7C+oBwh
aotoW+oVFfOUE3RtVsmydXZOYfCNyJ+k/qCiy1whnk+SfGrlYbIh/MGOntVohfqAgbAZNLhn6+K0
aXeHrhKCqUgm56MvpXu/udy8i3BNRa8x+phwwwsdA4pbv02czJXeK+ohFVMJSxET/kAt2/h3eQ1w
XC+tngmgUkNvi2uSvh29aen2B6X4n8hBuAZmVYA3idzmLiEzAAjBM0Z9xiSp10Ug2TPaR0kaSJOK
DEKsvPrVaZcAVuiBZZWRAVtV6WZOKTMPdLv4MFs5fSlh5f3wF69F4iP6gagwiOhSNlBEhTijKQpq
Jbw4Qax0btdy0LwkUgOiC3RW7SJ3PKKLoEZj26fKb4yMUqsHZRxJTK2vhhWSfJrOPGp65zpDc3zr
QUKLi8airUkUDWoVBeGea4o8L+8lPTteqfl3fHD3Kzmav0AIObiHhQV2g40xoqAonlwSbNZ3PTqG
Ll1wha5tR1a6j151UuA2AlOyMOM3sUZsLl1WjmF1/nhxR4pXaJe6CXFqKCsAgaRaLZ9tvs3uS4tj
V00Gx9ggsx5uJrVa8H7tgirs1czlajghR5DK7+OFahrgdg//ZR/SzkAHXUpFAluB4rmYHd/t3O7M
fFaQetZ95en2InHcJbKseGhfp1swaPkIXlcJPgu2x7xTWiUeVn1mBb4pW+HVK0Tyq2q4mQT056Ww
0kvlUQwbp69g5aAYE7v8V2171zLeP/cSxmqtaTZJSnSY8YUCcpRVc0ZkinMdA5jG6isIhlrcaPMH
oewWCll+/0tWmpBsDUkOlAFmE1hFeod/+62dBUfZ2oV5pWHP6HB4iTtsRu2JXadwwJJalJh8hA6e
fN1IauFCsq/cAUn4PZHT0f2TaYozfZugQhH6n9gsvHpXBpuMGqb6G5OmYFgamphHTsXy6g3SFoaP
6aKZ9mDVinSFiSCIbYPhWvML9AWDLKvmMjwcZrIirGD+vzoJFwz2Vo3pmqh/vq8+b0v6ZzeHxJWs
l1HV456ZjWw25xHA7aSmfCyNqAD7ieClxIScKMnEgXzLJ2Os4waFL6XqbUXWFeWiZRZg8E10yJoD
rt9p7/Ookx/X6nrlAqOwNbSVgYWRRY4KKcPpsZr1flkCa21rAv15u50ysFyTgwvMcEl/D07/fWz1
b85MMuhAQfN9Kl/jpeyOMhLGcst1jd7X97pJhflqK48Kv2+fHliulukuDo4Hf7zCNttCdMCRHK2z
9TBPHqydg4JJmdfq74fSuAW5bk+iZU7/ZwIOepvTfQ1vzyaCQCeTb3BG5ICGtZlDGpyOrR0T0jh+
ZuwAtOFO8f0bkl/HrVLxYkIti1varjxSoForqzhAlah6HluBI4Z7tf6JUZeRRa1y1HcdZwHNWA3m
78+qZgA6YJeznLwi7Ih3cHkxPGpg/OcjASIWhPndCi9V2eNndKif+K2BcoNoFCDc7845r/f3yG8d
+DosbEz28sYD/TMTHJ9xLl+5vLs/5tEWrB7Zwx7ArYMh10yCzXWoLo7JfPk7WlZIQS3Ku2v+a9Ng
SYhW+kj0jkUvkAbc4esbCt+qyjTFO3hafiUhDrBixugOEEDvH+qWmGgArIsmCk9ZtVRpYzrkMAsR
vJDuEp2rMAWvwFaiGUbg8G7gJitN0C/6DutsxpyV+7XGlT1TvbxC8MXIPG8UOnNHlw5TIMHaL2dQ
ZlLIVSmOEED8axdGx0Ji5IPoFjxpZeJJIhpXQ8NxG1Zr5KTCn613vDtXenE0jsjaE4U17KdRj9Qo
ofKhcosXd7qltiJtZB3Ojjdu56q9It+5xHfusIBPoOAihJ/oauWwcoShJxLKYYp7fZK4/W7kl5b4
+qDqH2MIGBHzH/OD8POdZgyGNEVGftWE7pPI1R0GtHN6o8DG9XSJ8/zSH/XUn9Zw3YZ5uv6W6+YZ
2jaZ8KCeCbiQRgYssd/vYk1w+1vMskad/eJwa1O2gLQqVXehqHJXGsD/rm6M96b2lrJJuRl0vlzF
qlWOt1pA0oXjk8VNP5GTIdiw5tvZwhDw+7cKpokBnq3tTj6ApOZn+++jJWrx8yvmXJAklC0kwpK/
CkwlPa9r3V7ieJdkAgs/byFnEFoJPe4tA7ajZ+VrZhdn0KvWU7zVbSWET5zZ61oecfdheHPCChCh
Y/IZz6RPZ5uEo6JVJ6a7tAilbm+P6v7tB1FKwnKLiMR6OjAzd0wrsTT5hp9QDJD2WYlY/p3hKL9i
O/C0KNax4r2YVTcGqt+VYxS3qIAoVXsuwq12sZFyHLAHuQSqShoSJi9zgMTIJrhtHZPEMTlq4Rws
XsG8TrfzkKMU6T1KjUnM8gN3XpZQwyxjMob7tAet6WQwFrk9hsvFC+/khkKh9XCdSyW9IXc0MNZv
flQhLb9eOdiY0Sbv1ZAyJbeg37H0LD8x0Zc2WFYd/0fdG8bW208Rgps6DMr7hpg6+HW8Ql0Whl/Y
7+1WvWP5t1RLkvBMTA1zn68aUttbLN7IjWohx+gg/zTQiGL/One1aX/wWnWZwmJXGqbGPObkEBTY
elxJ/aLbQbFudcvG1bXYyUsUoSyXCJGfin46PDvOVEKLIL+iy7HXwRHHrQuXnz2KRCT1l6dcqnyH
og9sz19qrrehSscTU/L0c7SOPL4G7aoczd+nh1KD8QpLChPLxIQPObUfBeJTfjbwsPjWgvs3Qvak
lau1BkS+ShvO1DXDrIOFfzQYc6qWMzceawJ6uOqY2PfwvgAqZiXf1O+JPimK8W3sPwHCkhjFr+kG
dq+vB6Tg7w0AP4d+8zWrpQTXHcxRjMpkqa8eNtAPLpoP1BEtznK89gJebEVBPCpGF6/XLAimGf74
08tSyJcf/tPFws8iDD9+z/jq0xdwXzEq8LiR4CavtUQ9lQSQ0yas4sMZ9roBuyd0KKEMlG5d5DGk
fU3mfh9MOF0ybVcJGaFu4G1NMWEXzuIZMw+UK5kpClz07bwyuRjQdKRdceLiuY352ew1/YpEq4tv
o/eeMvoiT9FAQ/K+H+RRjdXqnWFW+Z0PJVHza8vViiuZbA66BrCiIVeub4uzG8VGoxFAcGN2lYDj
Q7rUyYEQCnx4IpoJQpZCPx4ZqnVQll8ERVK5bC6gAm48/JbHo9TNtiI6KHMcDaKK7CuBen4Q2+DY
WPLyy3aeL/aJJSSB3MO1YztXBGP46XUB82I27NzjHKd+o3i0efvy0MD70xRizJDeyNZjonb4Ejta
ZWvuGbVNajJ0utHLfDgET4HvT7g7KgRpl0zMmfPA+i75jHFlSa80Yd4X3ZYhJ8N4WOA4yTQymDAk
6Qx7xU/8fNcRBmt93+GAanHEZEtemLuQ07QjRt9gasQoCDooEVNprZnAokTMxFIcOxZgUQCw5iRb
QX5nUr2NJu2JpwyO9zuTAi/k6LGx3rSqeL7/m9u+KvqKibGLBisA80k/da33YQpGG664l2JXNmHL
VVOFwuIH6psbewPZu+Vdhliz2qp8rf4Nx0H/jaa8JNoZduhOMreN3pgJHJqcA/8MS71ahLQ6yIrw
LI9twhPK8uUWZ2/VEIbL7KcHuhbQ0J3U90kDBUuOHzcLxpPWWcPs5u6p8JmTuzsqe3pxKRKRYPoI
oyrgOTizXQogltN+4+vP6EGlJ1zEotqeuqdksMLIJZOqJ6+7KxiIO78mmJ8SVONMZ8kkmKeWJ44N
6YplEfIZ0sYvGHO9mQyNKung57EQGTyxHaCB0INMiVnzhyPU/5wTuJZdA2Pi2KdpHh+lREtOjYur
sN+tc+EWurgw7JkuElnw2D/Izy426hNaRtW5kFyRdBw66g+/HDVXLXZBXbFEK4xg217RXrrcIAus
mDPsFybpySzFLNsBXqqjDp7wnnwNFY7m7bHrjoxAGAMRYyXzQdDU9YTr1GP7qFpTTk4U0nT0tRKN
Rdnv8fZXMNTzYWwCIyYtcjQjyzW/pS/w/2uCjPdn46ynxXsMNpXjUypRuPhZkImGtYSL+2Z06aV7
znPv4d+1pRpz/7imqHMVqomlo4Y5L0UajRPXH5FCqfEJFwyQN+ZDKrespywxFafdaTcQeOxnykqg
BMrdoRPKbVGz6z3oAPkOUceI6icwdEK29rL6tp5Pms2v0BCFyDaQ2XxJ70BbkHPDoitIyxWXUX/h
kBEDwWCKUNSiuJJSRXYERVrX3VEJP3vr/Ed//RPI6bD3ejVayyZ9vLC8ZxOamuZjiR+AHqn9+Lkc
aJqj4gnDKqqnnR52swCqbXFZDytvFCTTzbwlyNbnPDRGzDDjC22C68Uedo60GNvrhEw6jTDY/56O
ZxLiYEu0x1GM6qwLjgRfybKssEAMJia3BLopGvfPU4eieebnSyiONTaOAvKtKbqBglw1ms69RUXz
9WNPJU7gdRtJSmEke2d56MBMXY3ryS6BOzcaKzygoxju0mKUZcJEwiHDx6SY18zi7OTpkHodPO36
3im0PCbGcemCumBoZmveOIjHC3CzKdki/kjBVdCbwGyYFu87gmYEulcWKOZZOsZCfDgj9qBa+klE
dXyUi/ObonYWtS2u0K4gqSaQhw9W9a+qkAWCWHm0dO6xe8Xss75reFzkTPpkTyEIr+xd8NYt4ShN
Yq++E0WRp28/7n43o8R9PdWZCmkMayD7lhepJDHLUUAkTJOVftE3Q6E2QBrRx5vvmph1ZWqAxUeG
zzXBJ/Pnt43fX2lb0apnUoVMlfhKZ/0ENvQ9Ywz2LhlgGqjfH9R/7kMvmKN/Cn/OTXb+zX6MgEPq
wqi8toBBw3lLu+AiizeFWWevhLlLCeH3xW38dfemFV9Sn6HpWyi9DsvNixiNcQ1yy5LJVJhSQhcJ
XPJO0KrI4uvE4gP3tqsrCzGwhq1ZAGF0aHbyGl1LZUZOb6flwTK3d8RS8U/cbCGAZgRi79R2Wq0a
ubxzdAtExYu3ROemamsZJvOGA3I7NwgQm68atGZboRlDqLo1BYBv26NPIK6MP7OxqgQlnUve3RZ/
3hKV9slKx84gXGWgJcUWwPQb5L+KIdyqNK9aHiLN8fWeVwPeI80fPM7P7UIEswImzWfPegF2BMRm
0DT5h06e0Yil+66HjjUCXTv2/0PwjaMez/r1GwbocglfUTFS/O02BgPwiMC+69fIYcgJ962AzX6x
GbZ7ZLb0IWXatSHtKRJFz6vvPMq2RLo6ZeiI7ZWIvCEAN7yDdC1XVP87dOPtV3eELCKXwwt0Qg39
pKChVkk1b411qN3/g+6CSh03GXFqdZIuTmo/K/zCrTlHbfB2jSIYPQ8PGve0f7GzkMiwUbt+XHQp
BeYurVe9eHfez5nvXGZs5VGr47YYnQfbQO+Aa7xRSXUPgWJOFPas0ajqhtvGN2gGn0eT5unUFZ2h
4TdwCRTVg/rdtlDHVIpLfLlC+R4HAgp7w2KFXg7rJBF+eUYBNt9urA0OD0X6kb6bUcqEphAnJzDu
T5EgjuSYm7R6PZ9on/VZooDVFicl74WNJF06nYc2faGWEySwr8j+ErnHzrP/9u5/zYAjbmgdZqZr
H4gxVI1a4ZhfCem6ac1OGQd+xvSt1ojjYj0aNX7T6e9u0aD9PoxrbtNfA2I84VCsHz3ZHv5bCqft
hJYSLB6sCWNxRbWqFW82dC+0MQVxGDygBoh6BIkHNJxjZwla7uNtln5yudgQq7E+6UvftLtV1lww
jhKvtRghhjuEVRdBV7AQ3ZsgKvXOLIGuZ9TqZ61bCa+O/znaZztAKbuda7aAnV0GHKDvaHPzpG4n
zHT/VKwUffNA3DfwjrxWkP4zRMpmcFIxcmYLysjRicSx0dDn0cy/T2PdNBiDgJoxyfOXJTrzVdSi
Uaj5SAToYQ5t16ybr8txN1eIYkp5vNNHJypfui8o+G3XJzJwaNsNqHOx46T5XB1tgel0xx+L4WRi
mSxbvsqvBR0t/+AG0rEWhalezPvkOehygg61/DhiznuO1RbFa18M38IdrmwR8+7yXz/WZfguEl4D
wrohj6bM3AfAJ2tOj+tup9ENZvzK0WOU2kyxP15naeXd/uuoyypYPQG5Up0ztBADjP1NMutlXsja
Nz1UhSTfTWyWjLF39ms2CcFyCmgXtH5ynu649J8DbGGxIeRdp4RaUZkXhLM2oJxQgrCozh65L8+x
8TWp2fyJPLWUX7kJNS984p2EGfUTd2bFcH+kYns/tfEcsvWjJT+HSO2txpEIW4DMDUVOUNzOKWLI
2UmKoCY/AFedEf63mQSN90S5lnJRgCdIRl6g/Wd+ZGmIbOUTe6hrltMqGpimC1r+ypbyHIcE+GSi
LSbRlp2ePHiv88ItHfC6PGbgPiSSMJvde7+PhpxQrt6ya6C/w/Q4QDqUMfQVaDpyCTIr3yUWPj0x
yPHFE/RjssTMt4hX1Bg7SQrCxIm6D9vdiCpamQwiTI6BErXpM+nS3Mia0mrknq55RJBE5WZoTEuD
6fXFPeBW/ulwVVSmDDSvNPqqWXfqaHuNu4dfDJQgMcnvDmANrgGIvkuWQ76/bQO6lHdruC89qcUg
1C4WmVM+Mo1Cb8+Q9+UnMOCvLCRhuaGfOuk9b8ED4A8E1pI0CELPfqAUPk7FRBvCb5hea9aCl7N4
u/XgKlV8YKPf2fxP9eiuOOVN4ZbUP49lKbls+e01NuoRPCdDPsjG7BGfwuIYID537FrPJiq2wQGh
7DCmYnSGjqNiAIuSO5+u+qprd5yte3w8OCIBR/7rnto1XtUpgrXZ+GhFBxLiE/lRZvESN8ju7fuN
boN1MlzrT2fX+B+hlU4n3lR2dc3UM3ZP/8qgb+MEi315dtHcrZVKaGy/v2Hr7/dMGUB+DtIoqxa5
jMXRAnsYofnxYqsRekk8p7GlMfqTrifxByBMxKGh8gNBrMCHkDusF30is/BSvvybNlBhCObVtk/7
rE1irHHDbQVlFzYLyt2RuD+jwkyvwD7Nnl9ifgezH8/7RdQshdV2wwurRc6wfysjZ+W0mgWao3HC
LWt46Q/ypHrMvl4fkBKzA6HWPb/D77IcQN1h1CZqHR2W1IWrU34c//gR44+IxJsapY0FisNlyGSc
r9/zU4G5LDNhLdwfmKF+IXmJTg1Z/TOAdgBAOTaJfhJD27iigqwlr+Bv1HpEzdiHAlDxniJ5tPxK
HqdoYVvNUhj8A+1/Y/9hQ/qp4K1q/5akh+Q6Y9whu9tsnxG2Gk9VGoXRtURBktfknQ2hXhnIiSIo
Imue4h1Js/Rv7Ab+jT6MATuhg1dWShELmuHHcvBMDoHelRU9oC2b/T+UDYKgUHmITYPzGdXChz7a
jF8QOvm8N9BuTaZSBw64xwsaYHfdD8vg+fkb2ZM1tQJbhyHOV1duDtx7J7t2UaiIDSoek03SgDCc
kld1sMU4qcsWYaBy6MsRMPBq9c7N6K8CEwIAEfdZJ6IMaN4JvCWzgR/M0Ahn5JkIufdL9g2Ecne2
rMTJUFhPJUMkq9tJunFBXu5y0M94rzu8X2pmg+iwvmyksxZVp1Gy2Uff0MIZc0ypRwLxlLc9v4Cz
P1DczqnK3zo5KfBoYqPaGBxSHaKhEH+0oIekkWaJH+7YIQwSgkjbB1Ei1NQIezqHVlAv0pEZdt4g
0UHn2YtQXjkylOjWD0sxC9SNBzLNZ9vIqdnMRTaQLJ3+f8KItRTHsAKo/3ZspfkpZCteuzOxoq2C
VaKtySTbjJahQCuBc6GmMIF9pXXTSMfKNZO3+I0twj59Rj17yg5R5J6kUrpEMAAdDEk5OD4zTjeK
+JtyfnKR4ZMxFOCr2C29d34D+PoDOLPt1x0gt2ardM/G+Qi8ri5ZGkONata7GcI9aEQH4XpSqyIY
n+mr4eryT70tQE8Xjy2ZuFcFQE8+bknaGA6gQe6wkRVGMGl0e0Im8R5vkLZ1G1HWBDLzIniFuYjv
o/3L/5SRhxUDF5vnSIf/Nlb83/1PFeY7xYjhYVGw0x2nBkuBxU6iDJNTPyzXJWUVlVdnNUnXqX8t
EqNQuib6gc5kaUu3y79AC9EI2wEf2qKjmWWGwNKVR7RRgcagYKZWtpIZFDZBwieggc2uupaVl748
TGEJtBqnFG/LtPWnCZjbIi3iuPCKG+qo7mWdKEk3kIcQm8De3Udp+gfGEk9Z5vSi0O9vKb2wmoOG
sQZ8+mq7yautOVTrlvdACprY/gVKhNL/oUBONCxEmQllL7rwegG2r8sbRiOhcZoVZhIeyzapWrpX
QQO7r994m0ieZQ9WA5WKxaEDNdeErhUCeYl+LBrVHaa2s+Q6rXngdsAqsxuVq7VZONELVrXQJ+sg
huDGe7gzIRqPbiiUuFZhr0/8YvT+durKWUT56oXHPj1+LF/AOyB7bFgvCJ8tDFOkgQpXXWZtbQ3n
lw0H3TjM1SfsKxXz9j2c+y3Nf5zj8X08iTkkt7wqM2VeWZJ0ngaRkcD1B3QCuDCRjPHb3IXWrWmY
M7AkXyFEEo5snpyGtAcIPkaBuG8WCEWplBX277/QcJ6pXj7iCnrVUfr2iCITIeUI/YWujbRl0kZt
UXiY9/UctFA08d7sm6+8sZeQaI5rhN41zdGTAGYjoWwT+NCPjCPtDrDGcs+/kBaO2cn7Txtf+abt
BY9BsVPqaf1haqWpzSA/VoUmgpm/qznHky4G2F6VIYrZpvgRIxHLhE1SGLrizq5qrBYNKjTMDU4w
FrS447IoyaWhXiKkyQXAVPrBvfFPkSZZNKo4k2POMPi/smrCTFbUxD6KWHBFwlsFjTNB+vJjIGHs
E2hql21kz6jDp1mGQ1ItGLSDAPzVqKfpbdSpn1awMPGSlt2mUJLeHjCjg60izcqfcCXaQKrqn0i1
HMnt608FU4seUoPAz8vwZSg5+TZYCx86uoOa07F8OUfx2d8ateMdDxaHykl8YKXhWMFJWDztk1CJ
ye66faBwD+d0PNZXCA/mjUV75tioLYm+KypvOEqd4DbK3DY9wJSDVDfx9feo5774mwn+9gcB7L5c
Km9jiLXUiHNyDBs5tFfdGJaUENO9NtP5CkXJVAo1ZlCqqw/GOTIPaDuspjg82ACDmND/7+eB9/pA
6Af4+bx425GOYSyU3qpInQVtpTeSQTn7b4Juz+ufdGTFHgNJMjWYgKJLnxDZX7u7K97frFmcaz7v
c4airrqJH88JHe70t9Bm7pzqMQUgHSjirpDepTa2ufK/ylTP1LF8DaARk77vuoSZwuHj43FVrsNJ
zkDHZGleOfiQdjJ7bKnueWd1bQdn/hop435jV4g1bMNjRahElKhegQNiFrF2HVrMOXowmbshhk6w
AaZU4Hz8eYjwNVlSiK86YZZz4ZBcGsC+fPjboKVe5U00wMhakq7C6AsALtHJxxPU1nMGwibB343+
MKicHAiPuGe1y1wCaI4Ugw3J8Ktnet8ZPORn+E2Hc//Vm1JpOcpulQPibI30MiYwyT6ZMrL951VE
dNLx3r137h14JfVLdC5FW5YfjAb5izwoxlxQx0iu4vDEoo7xLcFYGmlHZCob07scj4bo1zyvJGK7
kcLQvJT2kZMQN94zPGDoxIFZaqNa/scaBK6cUex82+TIKrgHycdDBB1ogPXsbYXS4mQyuWDsH/hw
7P2oWqlAbPu6ltGXqggFz74YCoH7sJ3b
`protect end_protected
