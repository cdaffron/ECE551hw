`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Cv28uy8joE66iuPQZmynXGT/eNO3zm9gZ6qfk53yyDqU+cBPaWBGRalDpEl6ipV7IrsrYAhVt4dm
UDqZV9Bbog==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a6VehEIxvyopryQ/lU+/MPou+40hUudIzhIEDAVCfL5Ia7qRt7XvdEX0HoUxCj86KTbBHdpOfevL
U5P/VJePWRjVS9SGOUffxj3+OeM7iXwds/2FUdVPE1UbTyKT8t5Lk178Jr6o7WgKcY1UBugQSeh9
a+0obOylm+37diODF6o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QsvdxbbjTUqIriTWaTw6B/gO3sW5C+ekoIJmTHUvjuCZ/VfFelMsaLwB2IA2fr6Oaode0MLig6vj
ZXktb+2DQGt7ZCCDPQ0qMQ9tF8dj05nhe4SaBu3rM96ao8RaoLFg2VpRf/g4mDZRKN7JPfvnIuox
d7NQITqfRppzHILszA4jTcnkvRGFEVnicbLLzCOled694TtFDm7bDVUWXcCM5JNMYly99XQXY6Ei
qCy+l21UT3LUBj4LxszY/oIERVkJGV+kMc08KkSYpd4mWTaP88Zd5v9I5DS7BZSQL5b1nNtS13tf
VVXzgQeVvZC30z8ij8mN4Ot2hGmP+wEIwpF/Jg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cY4uUz9I//T4yoss6dta0HQf0yl5duGhYmVvXqXmmwiBwkeh3PsWE0TZoWyWVUepmL9X0bG5+YGj
3celne7tFqeIzZDFw0liDFu7+MEkiTNrHNtc7fnEv9jcY4IDoub+T4CXxiXQRIUyoFZKyjlhhEHK
oA0nsG85+nUcq5/mmS0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BMebL8YLQQILEjHSjM7S4WwQckhaxutyflDuEe80EVGCU0omHWnl+vgrmlxLC7iNctj372khQ0ri
Phz3DxmGIqKDP2xp/rzcnMSDv+hoUNM9poxEJXT5q7f00IaIU5wpKBSQzf8f3OAtuf1qDDxxwbl+
lalmmiekWdYni2eGXDbIgZjUfVYMGzDlU1UPFVCOavA1crcKauYnVrJzWFCSN2BgyA7PkJ8B1xia
GoefWXm5FvJX2xIZRwecIj1VC5BmUIbMks0SBLSK/Bgj7nPrUeR/YNwusjqG4wj8TIvwtyb/Wdfp
srllk1eWn/H3x3mNG1fNwxrBiQ+Oe3MXnP42rw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59584)
`protect data_block
pnZ/77hXlSM3eVpRHb3a+SJVAcgjesur6bqQWqC54H9Dphz8GnpZLoRyaQq1ioIb4Xt6Fv4zooQu
x/NR5pLT+/w6pJLOiMT2ysRJylCxjME5JHtsi+awaqRlpQjR5x35InjAImFAzOBfb8KPtwGzlE5n
hnrYPsmQ1m5PzBceCzozgb2dPro+tntqvGWl3ATSeC4WCBJJZGMDNIBXQDEQyQYzMgGjuwYdlc+M
MrdMjf0WGgi8ZVZjpTgCXQ8aUyZ6pHoCEkxK1dIU3LWF5rAt7ExDJxnx8/bNeECaZvqq8B7QX1yK
OQV9JNoo1gitrv9xWYzBwh3frHNbLMEy1fGpDuz8QbLfDjF17l3nDjtwDrKMGjIM/HvLcWAvqY+S
lwu8JKvSpsmskdGccJUqg+NE4PtTsW9WtPBAdSkwkrMvUnCOdsUsG6vW/FAVwYaBr2NWTQFQ5EWt
lxWDUDNW049SGp97wguOkjPLubNbBce6XcCFCvBL377UWuNJBUv9GZ0xodWRDn2BsZZTY3sTtQ4H
SZFda+25g+u53SC0p0XCZJ9PqmRg27ZI/WseNmkKyW1uuNsexEzxWVKfQMIIGCTSH1I++CZZhne9
aauqcXy9fTxHOj4I3iwAso5ZWpY79VU9iuteuGzAYQ47BdcBKRBE6HJZPiENy4fH9IQ07ZwBkoIi
BYKQnot+sTmyRgN60u7KamuPQwrQgi4i0ogazJdTuVuRuSSozuLrugPAzwyTtId4XVEhMqAX/pCd
XJho/D/8BzPVauwjXH2zBVm9Himu+LfS2Goec8l8eA8Gny8VO/uvYbokN0HE+7hg490DvHnDFqu6
0naOjF6WJqXWY/voreFTaU+bJe4RNOIcUNjAqzsI5KjPvRMHEWsz6HlAkZtWvGBiIm3FOA7mFEw6
mMWdRfrBG5+9jfdAcwWcoIgy9jz1CJwcO8zAxMiGXuVAThmfrxLyz1dcIcVAmulhjGyNMfNXXyC3
PLyWGCegchrOosIQZGWJ7lGjJHGfW6rNvTZJGT4ebMRN45eohFBXzsWidCjC4ksDpjJuBI1HM9Pr
MiHO9Dg/NRqwsrfBHvT/pnoAMn7R844l3fvFojCntFgAtiHWgYobdpt2/s61Ml8Rfvek1DkZuqws
HH4NzALjh01MM+J/VOq1US3UDx+0cgvCH8HUl/kM35UPnoKAohX51teUgJxB3cOQsIwyJXiJsIGQ
dq/reQN0wG9nz38JJGsPMW58I/BFsrpG1ZAP3XWRnv4OJWDrhR8tSLWFaQVqGB3RY7ufhsbqmZVR
+2q2Rpk8w+lRuVDzJSuj+H6EDFymBTZ8V8kk7W2h+XNda8BlvwKttwLyNDVS/1ETB2vaKSjdVlnY
3PYbkFBz7XjRgkxiOn1G0gomnJ1Vz3kFs1wT4AaroyxvMMOkQRIntqu7CgcfUY19JCNig01ygv3g
Q3YA8Fm3U/KYI9tfrKtkAQkZ0gJj2TeNL3wI43jRe1XhTmkeo0M+RZGSZ+NbRCEGp0OxUyrXVU3p
yrrEA9AivQs6qDhhHz6D0SX8gi9zRLNqXXnMPT9hh1uMN+8v6nEocpGTMaGUM5d2XtuwfEes4PFk
eYdsiJJtr/baGjqW7N3iKrch1Ws9GgZvXPLtzlCpexoUbamp9bqQLuqRWtuvP18vdj5oSTXVn6rj
bXHjp4YXVhk8aaOep4iTDJsvtxwgysJltDxAQS4zbmStT8H/YTY6uX2qhhB6iIoCCYAdW/9aoH88
Gosl6xyXL3ZVUMneodZdo+y42ZqCaoX6Wy4hFqYi5b4RQOjXcMQUGKipIbBgX4k9rxZ4oBdEkY/v
ZSwX3G9yMt5Fz02WX+xxc9ceL73wSc85Eush7yXXfZcUo48Lx+B8ZSpeXDvIesYZN2ydQfY4OCj1
ppRr1eYkuAkeO7R3/yh9f58aKOGVFqvGcTvnISiJZfuetvWwoIpFYBXZgWGMINGUYt43qEiXxYv5
ht4rFnxhPUKFDuZsXsqvo9LLJDm6TVt9RgykpeyTBYmU2Z9tUkOoS4UjN8nZRWDrpOcYjEkR4eM6
hTCPnth54edonidSHfD+aJccbsgLCd33at/QTqXGwLWGqEmC5Wj3Ox4OWpttrdof+34qIk+yOSna
EbX3wC8atScLAbjZBUeQpzEMYxmZAvZviQ8g9C9hkJz+nDD5msZLJjyFkEU3EUXOAdAjFJ6HH36X
7Q1R3go2QS03hOsbFeQCAGRZWnDBq8Lx6YMd4H/AzOdh/9ERJlRY7V6ua+XA3+ozmlB0g20e+cwV
8/ckQvue7R/018wkO6um9N+REAWJT6AQDT1W2/x/C5hPfPrau+wqnlIxPQn+HctK52pIiZLX6spz
2/CHYujE/btABhEdYCG6psc11N6a3R5kUAUYcFxk/yJzJSeCMKQNuAY0zgBZsjnO4QK3qUtSZ6rL
UOgQBdiYj+H909D4NrSMYEd/aGEGBCXzPlFr6z7lDFqQAQnbpm6KxOymHJtZhjA5wXrSaXFFtRfR
l2D9HKs2xS8nf5JsfNdHk8T3JoXpX1GQYwfTmECMV3r0rUH6SObHNIHP+yKr32BqWua0mAb2uG2z
zKZLzEYivUTfdFwF3/exTNmLd6TxRZO9r5YVFlUPWuFFCwMSs7ahlcY5A+hohXkMN86yZVZlZazh
HUAxOCvy3X6iUXyTycoW9CbW3cNsNqL+XoX8hPFj0vbCJRvbzt9ut90OzIXtDxj0+8vIHuxi/pXm
R7S675awIv52IVAk5kXSkX2jKRAT/FqwXf6S1Y75fScSAlq4bw0A1Q5jHcHGZ7nw4F1vqQAIeR/0
2+vdCHrytaLB+uyBRr7PrYiLReuIdeqPteA0TsV8NeCpOBClXcdPd3LS6x9m9ZIKOofdgCP0w3jm
8vX0a+8TZisPonzYl52HqxoKqb2OcoUfkEvx9KYIxIf4n/84R+dpmg4TsYrsEc0LAXIT0D6v2wH3
1J3zFoaR1rYFHKKalK7I+9raVHpUMGl3Xt9CklwQrjjLwrVESMiFqYZfhpQhRAVpQmUZHuQ5WNvG
v/645yKNwwqrvRBQr6gqg3QyAN6Sbgh67yZt6M1C+wpahuh/yp/OQyeT/l36yEV6LbFKywO43RN3
LPgSsH8V/ZZSAvlxhkwuyRHkEcUkVq1yIkk3tQnhEFzDtng0gxRRGu/659P8rKhZwWlZ7tQSumTh
uaLq/HmKoXCwZ3mMSIaAsYhY/1gd3Ufa/cDB7y+LuEpt8SME55sE5/6yLTG+/ffYcLy0KTOtsywm
pliaTDe/B6E55MXH0rDB0UaUp2oBgs/JKoSrW+u3iGkgNSGxCo6CVTSKAlCFvJ9xOIlVtMJOHzkW
orvC/EYA2bzOSGMSGQp0Z+X3d/95ey4Qc15b1rrdsadSp/k3P95n06/l+K3yDbfDX9WFreCVb/fJ
6Hp6EZ9xWYrcMczfoRq75PIC1dtPMO54eOy6gVOm0mos6ftAqYvA+jkER4JjaMLVMxs5vsDTKtYv
+oHiV8uh88P7EN5bdBWSYGeVKUcCNjWEPt+gQHmMHcd1Fi25A/NLJFj2UI+5qabdVvtZ23UIGBrP
+tY6+68W9tlPFOh66UoNMXUVgX1OtnMebWVpIInFQql0SAEvCrhsU7F7mGTdgSOvPRSzFuOV4dCv
5UvAPBSwH+4oY6fHQqXXe/KH3+C96g9rf+1O3vJQX6GYqfifNREe8Qm1kjZCTSSr1TfZC1EBzpP5
DfzLs2GBnDr0NBFThMv/06jJHv6stBqUDNOg+/NtM/kJJcKCuWHqoiM57t8BEJP0D29WSylX/8ZH
pzA0LR01vs6RhiZvQj1cAvFmSGIRDe7R9fg7tIc3hUYSAX7rpwNvDxOiU/SgIfi74zyXCMdTLDJh
sdkYIicyPe4a3kdmwgN+KFyRz0ce2bvhFcqHET3nG9ruXHb9jpM7Jctwr17x3jGRruoSHW7AFLi5
56W/1zYGe0ByYImw4w84Soif0Q3LpvdJl9gv+pfaJDji1ak72WQC0i87JkCoY0SrHPWNkOXRWxFJ
QlEsHtmtZAgJRpyTtIQzuAlgmAq3gDv3tsmBB/iHPg1LgLpMnjXcC90ewlyuii6Q9mSrJ8xLd2gH
tgHn1U+8+ihmePI0LcWEkApkrakbgfR9Cue7hSMPMA+WcPANUxCuOFINZ8brmxNVIDdS+RrlEdxK
HzNl7y0bMDa0HMSsvKwTMVpuOF5XmRvf4o2uEo+j6JgxaZOyG3cF9NaOpIYxImI+iLKjmZS1OvQC
ncf4c1/arudjWTxZC/kHqOI9NCo86XmgTCekxYYp3SPQUFZVDsHsGeUpDuKYMmQdmeLe+8i1UfmP
Suqcs3wA9YfYbDr9h45f5grJFc70buH532jGwGB8mHnT4cfi4hVqZkRPHLJ/hL/8qamwDKvYybBh
shaKlMV++Wg6QR5TDq1xe5F8zua9yOCWigsNSjv+F6fS+EGCd7Hx0kes9apzRKuHvacks3bfRo97
su6Uuk91tz+ULAdxsy0WOBu44sEPeFatUntlpqXN18JUdnVucsydpou5mTjq/HWUgHbZ2DAe3VED
OMnRVs8ylALQQEPTnDFSzHOsxEHBDkyNHqjWKJxHYEPSOVzBHLmvXYY1Qzyyb6ik8ZbJb9fdKAor
UBdRkpgmTjf+Ukyga4ujQTGuKLI4jo79h9h089cgdpL3n6h+fDrWtLEwZZY8BuM/vZv1ZtQsQBkV
yr2zkvJdk1tJHuTL5jZyAHuUGhp4HmYXo77tuLQ9JcpgCv5JPD+buLxdNMKXx6YJLsPuFPSyBMJ5
UUwJkk/v40P46oBpfEJkKFggaFPbyjx12xgGdoxFxBrMo+9jh2kLrkqjgqFbtDTulQs9AkB1ZigY
Ts6GFG8m1FGzhjymWw5U3x87aJDZXHrtDlUIst/nwBI4SVKwIotXIBS8xs6bBAmqaELVrU3M80TI
z0N+CQELsmZvJHW7Z0YfgtX5cmjxF6K6A/lekC6/4/MO+1mZPn1Oza/btwQuvfe+rtOcsqMgS1V2
4mtPsNR2DHBMxJsQGA0t2AMg4df0uAbS0VthhA5aDFaDj59IMCDyYzd5Vmy98piBk3LXWmRncbXM
nwXy1AjeYA584XGylTbXlP1dLw1oOchreTNOms3dVTA9uVBhawqmHiuVB6XMfP1HRB0643uw2wdU
6YbkuLgWiN+tjZ3wZnjwQo9/GrHtrY8GxlHk0PHTu8pymeE8spZqG9JYz3IRn6AwrWSoocUtg1Hw
Gs9OuDITCZyRcWopTD1p2Cww6ZQ/D2Dl3XWXOJ0iudgCoVputX3Uz9YTrEisi8WkusbWbHO2lpKA
nz9gCAfR30oaFl1AlZBA68Q7spWZ6XbJ+EOlyNKrPIgBzCYGBLB7ENBBZ5Rt4DjKaPq5jViYb0Xa
s/DofXK+yU7xiuTTKicIiKKVLp7YcNxkKHz12J5xfCcTkrwqKgZULiTcI5U9yxatye4K9FnA4J4F
1O4B1+LET5WxrH1zwn9J5ZgAzL1ruEB1JRZhkZwkiLSFNzEgRb/vRdqPRGHXSUgtKTagfN991t8z
1uP805DTwPcNT4HaIhTTDYVgoXszksckxnkYd4yjMbrtcwQiwdXcEJ/OKWY74TGMVXwM5EUiBlKQ
y2dlwJMcWCx53z5WQeCW7+DIjUnQy83CrEap2AKZpNfXJccvurWKczXfTrwFuSI48eB/hSpRk8RZ
1Ln++v5JM9rwI2lTICpOK8jUsO0cyKJMNvTeAd/UvgxB/y9nov51Ebzb51T/Td/f4r01jzTVcBct
dCHHyHhseIgiJicpGsRUQ+yHoSbU1hut/lyrUaADNTs0LdD0vGBJeD+Q2zXnhXqh7PmFKktkTbX9
yI6emWsbRwT8D1DBj+9FBYTew5SIfIx3IWLofcZ0x1rz7EHCeRDKpZFCx8nE+cGw2MF7veCx2sYp
dk8MUVqiSt64W+CPZuNcarM49YBnGLhoRVDCYJrdXuoi5A1FlZtmmsnnBsMQmVooxk0ybwAi9UxT
QrE4voxSZBSXbTNme6RDJNyusWKhxIjKw44ngq8PLa68rWDgkHWaMG3cPTjKuIYHzJ7OM9exmva/
PeeSqGCAo8dmdGnO8Pvk1NPoFpaJNHQhOlFXh8uyZco4ASA2kwh9AmzJzWCH3KHXltTSV2RoGZPd
v6dv4ANqzOwiriJN4HQxEpWcgZdgawjWs6eXNiYfQbVgvbpP6sy6G51vhqS5gThrRIsya/W9iJ2t
YBZN/3qGZN+X9McuaDixOls5AwXpBs6qceCBtLUYnYx4O/Nhpr6gvRrpx2vZGonp5/l0fe1KFNbY
3IQxQDsQxvB4yI8IEqPAXUdhgw8IcdZvQLgcJBaahom9A2lbfpo0wC/9wfHtmJaYtNAIuAk62aTX
spvohLea4Jn6dKxt5oqdsQr+bjELzh0+UiveJq6OLjZ1Og0w62npx6btPlSp0kTg8BUvp3uPztvb
hXANPTNysSuyprimHHJfaA73lHMlw8JvuYsvK8L6HEB8aMa77ngpUnzNvkM8v5PYpm8JtpdUp0Lo
Kkh7/8mdYOv2nRaH2YHQqTWI22LYI4oQcVjQBRDoIj1j2ZW9fmtGFgoJIxFo/itOiUYFwcQJS+4h
Gw5yKHvP/Q2FkrxxB1Wo4UY6jXOoD1sWxWDlqwXWn3THYsRYkkgf3cGT/rO6NS7SaVTlYInw5ie/
L20IwGRADqo81wMhPB+FkTye+mbE/1GAGfjZ8e/cv8vtilBdbohOYdGSXxzVBLgg1U8xZo4a1lJd
e8tdLkPOhb3k0V5ifkKZNIyqDb1+TXfEaQIEahfxBjjF4e1fRaU0OhcE4+7l1ArwEGSC65JDR4Sh
tTN8o6Pgne9N++AAC8/qHm02WixrtpJJl3XTKw1Ve/K595qywcYOvS1x12W4dYO7srLwQ5pldcV9
oLeD0R4Qm864QAjoKqr1I81MFkUarLF9LzSbtC6+Lupu/mvbYKzJyKROWqqIuM0uCzjIgEDDeP3V
/6FL5pHyxUnHNVB/jRTsDh8yBp/wHpZ1UoXQW8BMkQ4B9jNPHZ9vE/A4nOlFUsVWEurOZBfXZjqD
aKEILAnnPI8vFk3BRgpYF0OF48Fs37COzLgVcIlFca7X76oiF2/k7NAJUIHbt6DvujW/sVB2KpG8
5vSYIV9SQfSBEDUcpNtuIFomHy/MfK2JB44cMvFbFQcCiVeirTiwhmgb23Dhmvh3yQvvJzCaFnqL
Pa9jrriQ9lIHn1JL/jZ4YSQRgK1ELBNk+iuOvY1AfNMSmrG7wBaX99rD8Ee/DnYMNsMi5ZzRqD2Z
9Lx6gPoHc8qhT8+1uA+xRjgNDSHLqhmnDEKpsXKbulJAu+JKFHzIA6jildm469xyrJtMP+qikD5Q
rqf+4pXbXig2S1rDwUKJmseCM4S8QO1SwI1hiUaj/gCESrvWyW6PnRhd2YMTNooxBjXpIXi60Rjf
Sbgb4YDcrSxXiJAjio+J03HKA6m6nqdIzTIodZcWMZlnQiSIH5r+Hn32uAUO76nIF2mFGlO8sHHF
gGfHUOFpzuQaG2BW/BnueraSr1vGtI8KKn7w5+rMb6mznf1odPSWQqG4X8ndLxTne6XktKiP7koD
MMwLgp4EymDBwFN8a0OIPmsH4r0r2lPBvByeCeQm3SX7ijF1nptzRpXOgfuNkDOWCi3qINkIrzIg
AypWeN7wCw/G8MWOVBglb4dwhi9ik4CR9BvDGbS8kDMQ7rL9HfDb+1wu1URN5O1SNqyV2cN6WGuK
CsQo56QkGRHfwHNqc9HhBj1H5tarlXBQ9lScANVVdmoNvp1f3J6tQH4QNSObIQc79ysPzuHxmPdm
WrrMAHPxuU7XZvgXrgWUJVvZF9YLMhqsTBgwYT6/PirNnBBYvYkLBA/6e42pWvTvgtchMFHy62oD
5yw8Brp6WCXJYGrYIr6eQWLd/16hcXAA32RDVGjii2pSGNkJXwBOiK0f2SWWRqaFxs67sZoADLbW
YbkvEOUqw0VGlxWPOEKirdJProa69lKrK2DH2lIHK8yckYjAzC380aFGfI7Mb256ipqAooNx8RvI
QdXCHtX6tX5h5lQxUzuoWrXkC6ey+wDbR+CiJb1jdViS1g3vq0TVjDOBGOaxQXs/2nmrS71Fc3zv
AeFam4XUEr56h5VQJ+vtk5iYH7q0fK8ukfGWKmMENAgNClJMCfQ8x5Pwxh6p6q9Iv764SGdQyAVt
Ot71IM/hVkmEo+STANsP7UmI0aAfX9yybmt+DoX9TJcItrwoBDy+nSWCZ0U3jLCAN90z1bnSY30J
+RKEC8bxXA2xwCoFIUMybXV0zBvU0noqPdf8cIXDiIqs9cnU/OcXfmdy/eB0lez6PPLnMTYukZpb
CIoG746QFfsza3dxO/EP53Od2yh2gD/y5RHNKMqOr5U8TywHpjmhENWvonfdKzABdlYh1oK3IK5U
GFkEp0m9Q6Z2yu4yen9wJGJuTWgYXz3r6xrG4fHF99jKicTxPxUMlNVwufMYmCw1IkoXBbf4CxwE
pDskhKxi3Mo9V24+4xW+0S5DAJ8xwr+miO73CK3+VgPxhKnv3gW9fLBGCfchU5zsJeRyZGcUtzj4
r4cMZIE3OgYbeeg+ikdHwzMUY6hL3sADGYtmtsG7IW1jXs88x5ZkhQ4AIxP5H1y/7IqxvOlh8kIZ
vxve/efTUJ8NelQI4Rtv2QNfYTmF2L4Vqe8bwr2GfbCBCrzjShTJ61YuQUXELeBpMjcMb4rlSp/9
SeQGCGZgSKbOjx2aJWWSvxX/XiLLY53YeTRgbyHvK2381OFYWAYjh2lZp+UcQ0eq+nxH+06KcdZD
xcUMm3Oe1dYUtsVaPho+9ZbDXAWSjGjFKZ9JBld8Gl8cSRdJPRBgOi6HVshTODlQ7sqLW/ffGNhF
JlEYeSueQj5pHZ/YHNRIUybiof6cy+eRl2tnxgz0ODNiyZuxJzq9dv9oGoiuDN1in9EPQr/5mT4G
7usPp9YKGGBCZ+eendlUwaK5Py8fDidbpYjcjRVDuwikrqsBQ/n4/irMGgVYQR5/5C/pCjIvzpi4
WBiv6vZ19Rsu/XqUdACc2BIGqoObiCXpd2ITjB59imINXOBjFxNXpE5WRMDYAHLmwTqxg+kdBRxP
ezOyXFQoCNCECvoqxQTqgsdVTLYRjmzs5Rm8kZ0ztjCoZDfpbvctB1xZHaUdyERXfKU3BqdnAz87
YNZFjvtqCVcOFe+zAOBKhyjxPF6lLkOClHyZmbM4yWtXyU1fBiJvBwIbGzwjVhG3s7BeZKaRsz9E
I3Zt96V3suPPBzcXV+R1s202gebuUw7kXTwIabIChMfezF1Z87MQGjFmCHcyA5ygIk5ghqE1S8kU
kwt9ipj/q55TxSIcDWfZeUqE8U+yfeMUomDSuvbXSwxtl6pWzphA+OU9+phSYLBDDCCnurdzKIpK
HLQ+TOEheTLuRc22FVPXgv+kReCJlDUu2LCjd0YMKjBwaFwOnpqosgOrdbgSBNy1PQ2xTnBlYipG
xvtH/CGIOzArPxKHNAYNBx8ub/iYYqnLa7OOg+uTrhZNfrVfqQrvE7WOQgBt/f3p+ocZleNsqNlS
iH19Nr2ANTnxWmicVEyS75yKe+vkimJSU6fG5wW0IvXjaBQO3bsQU1RyeEYlwOf2kSHEVre81Bxd
xXjqFljOfJKzDwKTViBur2S8WccLudJFES83M5OpyT+9zuHlQB5QLn859QlidTWUaMgN6/Yrh/q4
tKGlDfqeprhSF8IY9lKt1n8zucgUBZ7QdSyoDBgj7ZLYy/rzc4qeC4KvJFiozN7FvZBdig2U4H0l
Xpw1UwIApzT6QxXo5Rh2a/PhQvkms5Ywep6Gi7U2H56+bm82Xhjqn+spNpE6PbXY3oXeJ6UWnCep
ZDScVJF9LFtx/SYUDqbXDNz2M9SCHpWpbJy51vk7dAsYPsfKmICwYp+OYPt47boHbNNKUV8lXj4x
uJrdzUsjO6jYb1JjBMVdNUHRb9eNqJ3md1d3ALRWfxIaTcX/cBwqTQQe99RGOrF7vxA/zM4tSH9r
Gf3/ChpyFxwi62Hyispua+7RA4JDUHCTMNVZYAdMSSX7NdvD8rj5oz3gO4hGOAf6W8Mge1XhiKuj
LlmP3qKeZfxFW1UalaARdebiuSndeGC76ZjlvntLcCUGBUwbDa/Yfb5CxHAjyl7HwZhn8/C+LkOL
qEEmEjh0spyTouq2w8d/0Lu33sB+kWTH2GDr8gfu9ooB6FzC/ez6SOnbGUYvD0PfOl84r3GNdL5b
2h8GDMBhNXs8fHc+Z91KYJn1M4uvC3HBTmtjDuLrdnbSyptphO+ss7zfcg31zTUTYFQyoloSZsM1
fi2TJfSUYza8NwddFt8aV6o8ofsqEqkTFQ2dGEg9Ss/urBFYD7keFcU63ICqC8WsSqTAWSj531zr
ueihOBURUNNBaxRV5pboNLATPYSMgknDATwKa2HQAI/jDuYenGNYGQ7X1A4ZC/PcQuSQ6qtq7oSA
xzhn/lxKQJrptxLxhyMcTYuQE4/sE9YolyUpEAlfUpUDKyT4a2fWGJiO03PnrSXJNJMLAcBP5GEK
kj3yBpsfwSVGYgtStipb20EVeDX1ZxrjLbnK87ff+IjSzYeFacxjFlCRm8w2ZosEsbUk8Lxu+ED2
6haoFYxWPplL+cBS19CKjUFLzJDec4jCeFvgqa3fu2dA8MxTunj6S++VVfA6U5ExJtf5Vo1U4sap
xpp1xd+CiY8WOJm0IZIo/dQqlh0Ko/hPXtcpp3QXJMfYmYxQhwfXCX2ZGiEJ2kgOHDQt7SVbtGd3
w+hTDDxXgOglpY1wsZLXpsCgyH+rbZJz468cgloZKCct7XW/qUbqaXNZT62+L24gJBRYuXsd5A7f
e9nlbA+jzJ6YZkNB/8Kjt/5FxvhBNti+Mo6w5VLTxPVRg0fEiyROvWB6XVKXpED9j+Nmj6IxFqtF
XM+bSfoWp9khsfZUAT324LJz5DhRN6tk2Gkb0Gv727Vt70A2y504Yeh3aJpjuKWbu7rMeNpbAyox
baSANqY4ZqalNRajozfveZg6BkMqJXI0PQhI3En8p9qSzCA3UZy0oJjh8pnaMntBLEXt3XjEm3Kg
44AeuJiAJlb4q3oazSz0j9T7yZ3iUauvnwOulYAOBTVf8O6zXjRXxAz7+0xI0pVNkPK36g6Pypl7
lb6OMRoZfMWBl/oOu36L98IminmPiEeSAZxTstPkQ+ZspOe1SHMb4vTWNbSUwNS6/xJ6eGccpl3z
bE651rL8vb0eZC9TFI5PsbwE8MoY8d2uDtLYe41bat12sPBmgGg5NYk6tQmBFEGZz1Tr0MED9/o+
xW18QM8zoZYziFEQvlmaRkBHE/WqdBSlGRwNJFGp5OGcReh+1mnsDqWdb5aWmK7ZfdMvjoQ3AHge
iIibveP8ivPFqtVKcrz7q5kLuUgkEsV4wMK2hNzcgR5e7HjNRuaFmgSf7wFPgv+W7zGfSwlpnuPN
uaB/1q2rHPpDX9+ZJR4lySUev1FfBL3Dl95XoRiQRwDXa8c+f8168Zi4t8nOwuzIuB4nikIpeBkF
LHyvLckb0rT656A3aIbBjJfqlp4h9fTw/yB4c2yyyaQRXvS3dK7n+eoGbZCg4PPEDAscX7FZ9HSl
NzTM7tiDbZgR5O8eEQ4HUrsAGlhkgRyfk7h6LXSV0aD0aYxO/ISEXoIP84on4TPxTjKRCOYrYsRm
xK0tRSQ+SPa+46/XTdNtwx9pL5kpOpDK386l05B2PkqMQFsgNMRn7yNVfVJZUCBdVsgR1bk8J6ym
GFuUtGDYlLw48R1EsA19SOsgrE043T1CKh5iOA4xeF14p55CWE1C3eqtQNB1c2VqTOwhprpzrTie
Wqm+rGhNy1holsHnvBdF29W2gY8cTjqbHJTvkghkPnCK6I0ZBc1Gfg/imdk03fvZFjrLRrMSRpcl
EETVWLgJ5560kkyhjtkHP3gDWXwaMGy/u95azbZBFQgAAYk1w49E0I90edcmYqDLRpzCxJYgLwl2
vXizFe6N+LBvgON36Vkh9xqKHYuc21WXh6jTTWZseeevXK5bya4U557jcEiw6sPdzIBjs1PkR2wj
ZnZk+r4fJ3FzoV375441+0teEc8ke4k7GgDH107OAssNOq/3T4PJqqTH5eBPQ4a+tqT6jF4fp7Ad
+1bgi4pig1n3ASGplycJVkYQM9Iq9gXGY6FATY0UVDLMKFD38kby3n3VA6sBW27ObpU0WQupVQK3
eZi+pyVUlvkkQJVQykt1ezOmlqv7L7nxNhQmx70L3wbbeK/4IMaSuj1GeQrR+2caPCrrF+YHVC9L
ubiZwZDEeEILtoAhA3tj2ulHPqMEC/Z1hwgzW4nD7mnFZUEynrkRnNTO5MaMN0tL0tH+EFdIObxJ
9L0Pa9loou9V1T8y6izomIqbT4yj9aseEWHkT6OGkXHx8dkuHv92YSB9Tg4cLUylejRs1RYu01fG
Zwbsxg/whzQXUi5CE0bQMzRGU8NreXHMhxuKGue/hjV/9kItEfmPnb/fR1kD8IM3x1eVhD+FZQxH
4Cal416KJs+WsS1hqgCfDqpqfEcOrG7imfPAKuRY6kvo75H7THxJY1sYWL18QfNnfBw3V/qQakoM
a88g68mrxt0TxszxQdIYxLsNGAtKrwuqJ/VQkZI4uLGCzwskoV5MA5FSRicSI5dZbdNktN9pCP5D
cEsRVd67RQLZBfjbo5ddW1X0tcSaHy4/EvBtNnx5Xm9TwEqBQkNqlWmGfENXWXpMCaFjBtaV8bT3
AZe56sOFnYh7Ef7KsaGOwMINGqnZTTJcjvJ8X2CBjAZBnBQ9++gON/XKgazswNoPAo6ttR8lEXaD
tvuLsA6ZPhHwE6ec+N0MvuxDbpntHkwcGW29zQYtw2QKLFp36XXxnQ003SVEgBjvJkPgcldTU5FF
RUzMUTDWwtwQNKdnMbSd/yue6OtD4ZXio6hoOMbovKLvSyxcsQNJ2YFdXlzcAzBWgFrSscuUmLPx
gQJzjnnZlCKuwP1dsl2xujSkPi8/s0faC3pj+jQPy1RaQKLInUfXA2UI38aPkKxXrNYpqZ5p4fT1
sDFfKB9uPHdBS/Y8HLdX52JyKDJ8LiU1plSRtJHvVfqhqkkH2NSPGP2yTVZT93KNtBtrm30X56oC
jHsaWiuLHQFHwjALwBp8c7GT/lgY4MGTPiNuYeLIEXjCYHKL6Qp3GrwGPbl+ncbqV6YNROI7l4fL
YhLw/Yx9plfigHhSwNBM/5Wf1QgAWKgsAVeGRlmZuW8Aqw0jlEfEvlVLzmOGzR/zB8jG02rkKM1N
uM31MlY2h00d9jmoTr9LMoCYUAjuCE3FmaKHIkjnBi5hRHikDWapI5R0/qi6b/4azm046baa3qBv
AMenztsKwRXxOLQa12xpj8HfZta5UWFbWMQg7wt47LyVeDrGlOx5J3LY65Srr6ityIwnzKBp1A5I
69lGLdU7uHqqCc7Q53lWypimAj5qLdbGbYHAD8wLgwqvmIfasJA0CMlMIofcPqTIKLnYSdUrrIhL
v5g/Dl/ByJraHFrRy1n6TGH4EytAzkSzg0wbmz9cqSJodJfk7VesxTeoEiRJVNXZMu2uu25UzOhA
YvkCxSAp/OPNuhtSewatHDnSmAsK5dlTEqwHJ+jmkaBMWMXa14R2+YH6XVpJ4f7xFK17blcpmU88
RdLGM6T/Qixur7zdRgJw6YYSv7UDrgQBYsLUDwrUMekqwQwCviB4RVW90J6/6+sGOmid2ezM6EfC
Wpt8bHXYBnZ9J1ITR23/zMT541Z6jVt7AAbSHTm0SY6rkYTSMBLLt0udT1tWH3nlHwKx/bM/qZly
Rog+JI2nE1G+OAKQMUjES3X1gN5603AFLb9i0PKcgd6pHYp8gLhcPaLRPxwx22RlB7CUeGkX6Fsv
gISsBj/KdTbBbwt3vA9JXG7J2u2kmQOJEzS/ydOXT+4Vh3N77LSiBij4sbh0mP/glVSwCjMl6n1S
ZpzDYENAwikFsEIY/X0D0mqxEU+EXLQN2C1ZTxYap6CPJ2R/V6OQsbDji4RPIzg8J1H4jDaNtHT5
iyCcukzRWQAPLs50eMHkEX1cM489UDoVjM+1nQXA+UJh9QdBLtibf6xqy4DtHbRZ7/3XqkjvSPUX
v8Txg6BYiZB7owmPs8gXg5HGDSC6ctiDIM9DN1S/iq93BOmCQJ4pY4uDkNaew1C9OD8fLmQgS8o0
YHws+7Ixo4FA94RMFkux+sA2BaLWDt0v2cNGcjUQNKnfVnZJdX5oT1tr5szgCD8JyzqDRQ7JmImS
z21XzNzHFUbpTrXH7EZ+2Bb0o6Fr3RIOASJ7ggNKvz8ybJXvxAh5vn1Kgtt3TmHNTnC1/kwEwr7M
HpNvBRW7oExJa4Dg0ZVewtdbSuJPJUX1RiDzjc/Tj4c2eb6Aqk9AMlWAWPOLH74vFNPF+xTDr26O
sHAyBsP2mVnASqGL2mSnSl1EVkC/lEqEKFo6qEq4n2DRKO8v2UOC1rfD64SAKnlsa0psix6rdEK1
LEh2ZC3ucmv/e7sXStsQM0xeVLXEXm8yYgRjmdJQZWDQqAKux7R7cVjzUU19W1Xt2y286qooQFb8
L5IjaF596jfrPQ55fOEqFKymApe/r64JZK/tv4h+RyMupmNRKkRM3JXBgv8fmeZRfiGEh1tRHVRn
0aTHvy9XUvxedmLFh2YexyaEjwygCb+3zbFbxj4R6TAoFU1jgFRaACHSxDHsc3WRfBRZYiRzqnl1
EvDiUJG6M7nlQgL2E40WhlESgc/C2vfTC+qLtepJhdtk73R9jv9jQaHdctzrcFVc8eFZpLcnPxfb
+6stoLjpD1ja08upjniaV/QlX0crMlfTOo5Gb+8dP37M0WNTM/tJM0czv8Ib/NhcxMWrs/VtbBcz
Dr41pCHaS4SlptFfaayAvekm047zRakICNBKq2f92PmLGxmnU+zTT7YgkWePKLqq5+1Xb7XcPIFz
O8F7N+HU7wbrKHre7fwfVlP4hbnPWIS91G+gVc1C2nHGsfZNFcfBe0RytpWoe0V14eQ32mtuTg/w
Z2wirx2qj/79fRw5uHuxo9kcq1Gcxe6xlIPnU+B12lb303Jez8UI9fqjdxzgNv0RMng8qBAFwC7+
whs2WHeudjD0mzXFYqLqWJOL0jpTX6Knnt9IwrtIdsqI+/YKLKJk6t8YlWucKX988LmWszyv+ICW
/nGL3+rDT473dameBQbC6hk8OA3UKgzU4cLC+r38zshps3o1oKR3otbj4hxq8hrSfJBystHZoHu8
U5sEmOivocW1zFCyLO23JbSgmo0LRLNJjeHNWqYIJlYaRA9bf22uu7rt9oaKLh+dnWILHAcVo6Ka
c7tL8gT27k9729oiXWSoR7niUMBOomv6HMMqUr4aQrxiN4HQf8I8RQz5wVbzMXdKxEaLAOOsliWv
gNBSZBKWbjIdFk2U+j8qY8m732/06G+6TWg6P8QK/yKFu/JdYhP+mbm+ftm1ov+p7HPnGuXRi6v4
yZQ2emSEIU+xX6XFpubZpdryAZVoJUxh3ujRylhasHyVBd5drXj0gnVNRKuuziqmMvLRRH49If6i
2lPuU3H8jJkkAb6nbIr6GYBwEE3j5DeIArzgzvUKnMaa4hk71BPRqcbckTJLnSt/mA/3iKAmwrE0
rqtgZhM3g+XXiVrpK2syITT8/2qMviRm9wL4nDFxnI/c9HvV1fOs0vYpQ8A34C7+ukXDaNWSg0Xu
ALpmXxJsuTg844H5RCawlFOkMacEzyI1240C0xoA4EBZQEz73Z3hbBDNelEP3l6D4qjtlQVCwfYR
E03OlVJu/0BS3t2CVz7CW2snp/be4Y9eLC8hQMd/x4Faj3g4botfSYh46Jm+1a9ZfNSfZ7YO0N1f
E/eZHbaKzzCsv7pg3+PHK5fHdmOQTnDqtaWB3kGArBN9hqNsZ7wxUvGNpFRDdsEoOMIh9Yiu9FfH
NVKds8AVI/t1pR64faz7Q2Zuhfl8ukKOKr4E8EmTA/jz5L2hlUSgeK0D93WwHmMHGtHyLm3e185/
xk13VVwq8lujPjyJoimD6h4tx3cqmqrBPiCEBmuDwEaB2KHRsNvwGLvZhnmTPju3gloxq9pOL5aD
WD0UFOIOQQ11Xh7Xw5kHApioT/lJE93dPyC+IVrdCpbuMeix56vS4BwhInJ8Sei6dC5s1X0mL45D
NxTm+5OE1jrbFoIvK7xwun47O6rjJYsfaU8XbiijtZOFM6BQJTMByvvRgRsbeDKRNeXmZeWE6vj1
NPg2+8CJ732zpaHBfh8paJJgOUZ2VqjZ5fLy6tts9x9vbsoWHf+LDFPY5+G3BXSpO6hTZDykT5hq
0lq+TLuCTW0vvf/wpdhiYiX0VJeowsJQiDkhIeSDmTtvF7hpYaLyD4OMIvEb7E/JZqjwUIR64eXb
F51O0mWZkOM695iAaTm7tmCvHNlf36nTTVGAJgXABQIqsz9hYwEV31w1buwmi3Cd51yehyhAssSM
A02n1Oq7j9Aw3kKwdP9sRXIfbA1ueIvxMkYyBz4jqc7u7lSc7M7DF1UcYxCP6YZ4SebURgpWyDML
0LbuyvUDf4O/t0HMDkzV2oeYYrk8INWrwOQilKHEkSpv1QjY4t+iT4JNofm9tmJ1FfCyABmWrDtM
NevYtthtaAm2fkIzXeClfocYIm/kGaCocXkVS1jGMM7PX1uSklgZbeKWtjQcnXQ9T5qt5BArNP5+
h4eSsGR9Vh1ibF0fdtR4yIuHHucCm1jk3ApEs7Sk1hAlKVe4+otSVgmO9ztVlGt8s79RGC2jzdlF
vx4GdXmcH6nv9nvsFnQt81cHzISpETtptRnMGehLhZ7bs7ItLZVu1jTWjaKnPKtfdvypYMMzS3UZ
FN32vW6FqnjO26bxhRsG9GJhwFuaKgY1Bx8wMquj5Xmg6QdnpiIQUdnvWsvUJFnpXWqD6kj+bYg+
OowpOlFLlDHlMxAP9NMML/ubHyBYeNmiRSq3s+sWyUV7rl9Nd7oJ9pYV5dQXCY+ilJxdyvNiMRRF
YQBaVign0yqwfPUSd4AteRN0Rg8L+xZAmghJMGL0goTD5yzV7pV9m8155rOgOtoGSzi+qTRa8vf4
hzI0J6Bc6sS2N1N7EsTeVsPjj6A182Y2a3t8bdzXay4SCyIKogp/e4/aEl3ahiMyNekriNUDoWvJ
LszThuTQVaD0DboDPuj9bRom9aCtSU/QBQ48GXoPf0uThxqKcPyaf/kbXU8R8TpmxGLtNM5FkXC0
EJFnpUpReitxDVwZaJlbG9xi0bOjsyoS2acOEkMH638BaEEHZ2Xfk696DJcp8XZxd/bjSH6x1P98
+dPAPMLT+9NLr8gtGzYt7idVl4QMBHFAxC0Ut4ddnoiFn4aJgO+/HuuRsfBFz8gronSgRenxFF76
t4ZVJVk9WsbrdQ2pAsEAcxYtp8h+e9LF7M2i+qi8J961hHgFy9rPTnW2AJgNv4M27SywG9/+pOe2
5e2AU4Sc5LVXD9cg1ztcAlBhbRiSnPrQxcShdlr9W4My50Z42356Lc49CNEN8sawLjgMI4SZFDNv
IT1SqEwRhmgacLGRBOqhrLeRlWV8tD4TZgkG1dMKcqdTN86c+1QiqHZp6AZr61wG+6EtaN2SjNIY
HKt5xcxdTpWbTCC8iqY3daqhXiF4xZxZuYR6H94W9IAU3M5/IVHkWaCAot5q4OgdNPiFG1wht4Ir
RlcyDid6AZlPaBluZYpaSwCm1yxlNaOu0qyYJ/4/UbtNjFPeY7f1Zi9y0tpNTn3nxpLlg3ysQxw+
yUQt0pKMnlV+GdQWbrR+Vt3gxkbRqyIfJD5bxOMWqiJ5AHRHX8zcco3t1kxdh0Vp0G0K9kvvT5/t
JUKWB2cMa8ROgTCW+X6wcPOxwZCIsgz3QpQikGvTMDAk0w5gXwpFTzxp2W624wGvmAnHHW/XY0wF
8TwoNrqT4Zir6y0UsyCW0JTwj+tkwrhdJqqbJh1/8ikXE1mNVVW/xUA3n/t1Q3Sk/y+Pdp+d7Vz/
7pf9z/APvPPfJ/HF9u7orhMatmSkakT5wW7sSOW2BlLt6xS0nKgvpFGrmyg+aGCOz/Ge1iktuDvf
DfuDC4Mm5gykW5KEY1/jZH+Y32yRhv2NX1n3UvmUJYBVhhdpqyRBWylgAe1ziAHzXnqf6d2ggmen
fYdpWfLzRUF2Xiolwdv8ZuOMlku+ez9bQJH8MQoNR97uv6wAAAptioNGPdIHuSJcgFuqSB36pVrg
5LSz/QNOdZIE06q5R8Lk9gbGk26yEGeVPrHyp1pw9P4xFSTkY6KWO9EfyqXEr02KuK1QrqMgZsl0
gm0dp7ReO2Q4AMAwNFkB38ZfONEKo6jBI1TFpN0+s7zVQqplqgyswon/ux/liy9ikbwSQwJL2u3M
aXyFRoofa2ze77SmZFm014XkljL39N72zmXOMIpIhy0JPnC3zhiK3JdPVM5GbJUeYgpt+wA0Hynn
ogU0ZggpjQZQIGp/6Dgybt9Llyy4J9QyyOAM77F1ZL5JIQxnJkWkat1fi8ZdYj/lakiPL/buVxLE
xtamRir/Wm01EHAeRoTnt9pr1K0zMghHUY4V1OgfC3oYHA63wxeDO5rmYAqeHBKbk6ApWQQChF6Y
yOLYiEnfi/yuLFpVj7qS8GcCmxaKn1osw7zS7KFIyLhHpb6EsTHENB/V87JOAQGMRc4uRIBwqS3C
/NZ6eC9l0R2FkkyR5fz4HNktHZL19gzqyVLp7cmQIPEVk3getMIna3y8B+TTHyoBS/QyRntfd2UN
VBFaAoshtej3j/NMoj14SLJsTJg5VgU+KJ2fPoSv07k0+CmGceL+HS5KZ2LpuXnyfmpBud8RGdjF
NkCvyY/aReavo/nN0i9yf/F+uBziyLDtABxJPZgBaAV+5WtmauRaYOtmAVpWw1JVyIgdZI5AgBrx
Sv8U5wNIfHo2QgVvEompAddcuBKzDJSYH7EXPhJuPBMZZiQEgewuLtSNAhdou13ILcqmLVlPqhO7
spdrd9UusWt6PiVQ1VxWgjflyQ+HjDlHBVraAZU9F4hq/X0PVUwc3gOzr3Daz/i0H/Ml4iQV0V5r
iQDX43JpRNRvvJnsKEvPqNCzkOu+2Huzi1nsK7XNglVANi7jYHd9RnNKY4t0zlRtUGMcvG/EmXS1
ZaR+vYs7ANghIBvZQGJgsnzohJZuPfKfHoV9UvmNwUXMGTbD+tnV48R6l84ubk8fiLR5yAz7wKe3
FHBN8pRspisGyTwEyIegsqYgZHDY4ASpBugga3el8HOo8k0lahHCl7uBu/cmBOa3vXuwSNMonZJW
QFytH2N7qqq0faKlR9UmvICZnxU5PvLY0vO9NJocZCGs0Az5Gp1mj7Esz5nSoChuBXSJ7Jd9jI4Z
2Y7jY8tWEj41af6n/EIPHBBgp6qS2BGRJnC0qZDeX68byUlCHTzjfink2I/oQnCw0GG6oxYIetm1
IYnW0CBiXD3cFR5cvTOHMHvjcVNY7kqlWW9ymTSoW4CwLxPOFSu9vwEwCsORoHKfie0YIEv99ZpU
At8HUnnHqh2Pgm2cn3+jb69SGol/MqvY8wMKotdv4/dVqzpigBbiXpA2IKFkmUbhXLo/RDf2K3XW
gn+R4aZw7A9C1s+J6O7eiXECfM7e3Y3PFDmg+x0XrQJckgNFQjWQp7wiQb+Sg5fd5mzgUo1cCIS6
HO87C70C3zTKqemVxEpCrbZEe+nNUb0+4ncKvvlC7q/LKMu42J9wTd77D6z3jh+WG1xN8MNWbUwt
796cDGFOrXoNX8pUcQdWU3fhUtTR5A8yuJ8CrHXw/x1KKrMtFj+rF4aHprFTqXSIwDDNonppuMvz
Yo7E/m+6IA2T4IzEore9Kk6iBz0e//R/6TB+dLwPW4MU9g1E0oo36hdrmpKYGnKx04m9mXSdRP2d
w5Ki+akKNgVAKopf8w4utaFe/gpR+RD9E6xHhJ30+NPfQsDjIrr21BqJENB48+nEWFtUQWpUawAL
e8T5GAC1DGshFGKzhMWDZ3NB9G3olHZJN/IfXP2oKTsOvZRXUvqqq4Sog896AkIIi6fCzmOwcgid
r8SP6rDITpto1NYBoVryPx4+m05anqic4JO4w9a36Z4XoL22lV5+zJl3qFvxr1trBRqIn9dUhSyT
OYdYAisJfy3UOrjbkTHQemnfbStRm1wYAie84Zi56hhIPH9tlthSEinRlQm8ng7g6/D6K8Ez3c0L
ae3xthuS9/LOhfm/WvTdxselhnt6BJqRJyYgDApG0ACsO1rweM6DXnQLZNWAfiRTZYlZGf4eh+TG
09L2Zg4kyyfO9FiBjxmCBOWYKNbIcdmhsBCCoRlkJpeKG2VNUB2S4gOPqk70fUB1gE4sD2dVkBTo
Oul1tpVo2SZYUsN4pjxRBK+1h7olLZ9VhlOomfHAP0L9j5Wo2wR0WrG298n6HPSY+0w0PuR22beG
CCiH2WWqc95hnSDHU8hFvV/3464kOaoKLXbHceO6brBt/h68hF2cOiG3aYNqCdlob3Af2zILYVKi
QYKalVgjyctubAy1qymXcY0iMFcuH6KIBC9LK7Y13M3FZnx+YUDnoSyC6x2Hwqz1PDy6dgvT6OfT
2ZOdfmcpTuE4IW/9DAspEjS66/wpCi8FJLBxGXAXOsDyoraOZ94qbST3C5BKlVBRNX+YpFRcb2pt
p6wFF0IwM72A8ewQTZg+DYy3Um2IIl1V21jwNqhgfT4KnNT3w55deYXtzRzqe/musSGEVVqGzptJ
69+sO1z1Arl3351lKMMZVuaJEK3dZ2cgH38yoCHM4NcAxtFW7FIfrKqDdMCPdK3Acg+Lfu3Rr1Cy
JkdtmzyUCwy+fIjZplaf+dlzOcVtukMo9kwN5gZI5XEejK/Ql+aFMO48/wePEURrQb/g7XXePcHC
UmbrW2V3cKikuPbJcAjBCGbbRLUcqCxhsCi+eMUm8Nx2YNVnPJlpMUzttKmlSjegvlF3HtVaueq7
MO0z99iBBxc3BEGaPnLgs7vvpC/1ty8uJCROEXjx2q6/DvlRAjg7453cQgemfZ8K+gtQezdM6E5f
7833coeHrC7gFYm1Vmis4iQ8177HQQcZh1OxdadmNZu3vPOixHh7f2iz9XLt0r+5J8Z5B3sUpwl4
t+1hstkrpr+T9NdFQMZb/MHiXzY9rIKPo/PWwx82p0VkVzFKJKwQ4VhLk1/NOmDxL/FX6/AXMlLI
wdqNd7onvBHBOghiSTTv5+9epJ018Tqp4dLkqc6/lgObtutv7U/hxb9XuRDQhHrJEmvzUkHBt9ar
HE7V/mRQV3HD2PI7OuMfpkKJl+XCpKIJgptSkqvoxJKeFmSlb61ovSZ+HsYXcd4igzTEcLEfY7rz
oRia356cHEKxO8F89kVXTLfvZmEU6ca6qhvYv0x0nQiUHUBun/984C+gLNzKKVyG/9DdMBICkvHL
FzwOqUrHzAkOoiGgp6jknZRffbAjV3e1lis9v0Ji41BCPNHvmzLYEwiWaSODw4nhLvMMKignOvYq
umrl+3C41vY+RB8PjXNCXaBK+AqZQM+tMSIR7S+HdCt+DoTIo21Y0iFwbPZheQNfW01NQ2RS9bO7
V4pePEtOcIGUaaXypqGdDkekWsYfGSKRoVM6BLg2lX+WjmBBzVCWIk96N/pnS1IQVGJWq13qQCEc
9f2vyuUx26m0wMDtvys/cChCkeBd3sc1Uhi+bWpeOV0fslgQz7GwFjJhLvTDvxYeBXKroY0F5RoJ
OeMcHl7yeh06uaVvHk2xq7p8/0fcO3uOSFx5AB8P/pbYU+AJDqADDwkRJzyev9IRkt2dPuyiNnNF
4Dg7GIQgI9ziw7xVSZ5wPDF20q4EG7s0VkPHAtJSxjs/2HnaFF6Q+UlWy3rwvxaLjiBo3DTltY/0
+d13bHpJX29qCy/NcTVIpSEGxq0h1jiSqdMcvdnEu78q4XKr4LZixfzFq0VkLeDryK+pAHbh1Z3w
XP8aKVfzERV9Ya3tHDXnhjm8vkTzgMSMjLcRU1G/uJeOEMvzkdjywqwftKSjBsnnt8YIk4l37E7u
62ZaHhE6N/04+IPpZEQ9syAs8vEJPiakuux6GNhEiTWNZV2eJwRuU9qPn1CBoeb9vXX0oUCeVq5y
RjTi7/TSvEQ5dxVjdPO5qQhQtWSe0ftMSmfYG735v9smdCppRvR1qP/qnVT21eOCZvFw1XU852+R
1RQv7teyv/9qO+YhiQwr7B3RHheJ98Lj16djjRks64fzNEP8YyETeWuIhdLh+oA9zdvqJ0tLB6r5
mi6bGULD+FG6yDY0Wp2QD9BxPoI6OqNqIr//5WZrkTPfNtMQdfYdqelhJWmjvgpMJIeTMVcjqge7
PM54pmFTGMgq3ScD+bAJaK1fzFlZLPrwgJIcr+gyrvEOTUCnW7gNB6esL27TPwup70YdHK5L7qvd
DX3donnzCTTW1OGj7voVfEsUpX5PoXAJtnlu3xgBKAzlNKo+k0bfGNdQfWAYi8/hq+9L9Rhqzcfh
ojjc4cjz1zZ8eKY2Dp3yikJ3nlGeI9v33rFKOnvDWBPY2ExP7feTwhwCKVIZ28YecKS5ZM3S47nc
Nk6pGtFuB3aUpKHItnWIttWuLSU0PJcrcTu/d234t3QenL/tQNK6vcQtztqH1S5hyQMzCnOjxLHq
voeNoelnJ8NSWrIfl71x8GkTetmhJMizkIONULJlRs6fSdMyV7ir5rFAatQrJ8zHyNVnukGXXt2y
FMe1Ban+i+s/6qrYP2QM1Dc1hUS5HXAI71QTMWwxDfHySKGa+iY6hDYGCE6ebLgOSgovpX+aE7HB
RkAa2pWsbegN/fyS75BXL65Zv5FCtcYot6hhtM76pXJbRyUwLfcBhBF4f6u41mwtH9PFpf47zity
Qslt3aJWevSQAuQk7PgPeW/3jGCErXzCQPJcqzTNHwZNDxtXSmDtudH8oPy9dXY1elTrYuv4Uvyv
ZUtNYLQ6FsJ8H8z7X1hGva14zN9+SYPCYq2ildHZVy345PMq5df8V7XB5zgj0zs56llJvR/9rAim
dl+N6sE2Va9CHfYQ2b1gvg8IbxM6eqKp3pk/Jwt2ySdQHpEEXLM52eDzFTVU0U+5LLEYVr2RD7jQ
XJmtHvitEpIxEmdubtI6VwsYUyOkcjr5sztSQfSURgh8uIzGoLKOJcWDqgTGgz62GWbbQWSAR0K6
woHfrq5n1FVKfPZVFXKWDZbjvNUG+X8O5uI14DTTxVnduFlT0kHt4/7Y6KhZNegS+YvubyFMSii5
GMcOz6QsFyFIMf3IgR805OCzLwCqkoXk1BomCi4rrvkNjNNeDbrCD1lChj4873hJTienGhBRErWv
/5VlhrCycFvKj/U5rXwA2q70xw/qHWoPq0MhjcX3zX/7949pHrde4QuOx3aCO4zB8Z9HaJDZR+SK
hpPMUdOT0D9kSolL3V773FD6GQzFP27mTW/YDWsZhdb1ftM2C5XQhAqCE2It2ogrxov9INEYqlps
HJwLRh0R/Vo4eB4uaEzpDfsZCVbyy3J/E40XsQL2qi5Rfq+8KyXS5fjZZd0t8pajxxiIsNXA23YF
Y13kdwl5/XGa8amgF/7WIreCojH12QD/eMLtJcFNMrTe1bQc0jDCJl1KDtzZU5Qv7CmjMbtRd9DO
sWm9PWjLyQ5jb0zFFg985mZVVfjT/qzB01URxYHyqYh2N7LmVyKKo0tlDAKNide7VPPZwMAkY2NZ
b0U6VuptkRUCpRX39v4FxxBi70Nu5jS5qstDHCq1iFKeFIGm4ppCpqzE7HiciPunYDwQxNYtcULy
kRPVPVyVjaSflZdM/wDlZGt6kaJd/XCH7iazdgr0k0no/gXdgOKNDttsSND6Eqj8IbKN+pCuZcyp
obGBcWOaFIi1pfNnMvvpiL/fLmrLEtCNhabdtKrJc5RhzGeMEm0W8ebokZCc5hiHlse2lBiGjWNL
hg8FmdtT2+6duBxt2RR+DDl8s4PEnhSvEf3oG7N0IhCsXPUiDGwEEdQVHMuuKw76jNszfR1S3Eha
SjhZMFDzRg4FtVmtZJaCcbNg98JWQNSFU9Td1OF1Y9k65JHbgjFGW14YfD+kuJtCbT+xttQXcYCJ
+Qh6xzHgDW7nMp1vWr37Wyre9R1jugHlMsckmaehrt1UZRIRvwc2bDHJ17FMQ4esSdw9ucQiLZEQ
I2Mzr37+iKITSdXl/Owp4wobTevYDX2j/ne7OQExegC9N/gKEaHb87bM1NGZL5nNFRHGAg/2ag4L
wnLx+om1bChkVCEBKdHBH9FF1bfaPK1D7dhVNXnrPJbeo3zo8QHqRYp+E/xLU0bfAD/zKSLC6vfz
9u0BgVZyvRiqjDktCmTxCikzBwopUJdoGNy5cCuwNvtDmVqNouMuSn1RJeyM4+ZjoOgO789Rmbr4
tzQKZAKat/lDatiy57XvBGJ+dHIqOktT+bpsUNFbJu+9VTTDLbZC5FXZE6FPwqMf8CXxJyGZiyVC
KWi5f8fHSdRk3tjGyGCyjcETgS8oXvJvpMQzslzCKG+cey543A0oHzd6Ilc+I2JTyeFPxeIpeSua
YuPcCVLJ/GTQ9hK7Ge938oDlKl7b4YNoXf+67dkYJ5AFPMSGU26sb8qNC0XbSEI+SZ53AHviRk4M
yJVw0wQTAzX30YfPGp+Y83dRq7CngW1Ke05VhjTheAJwTLwEaUDcM6W2/72ko0f2dPgqxFSEq7WC
gQAoUr8OWsn16wKZbaqrLSjifirt6DSNdCMzSU+4V+RMGdL7Qp4Qe+sBCcVFMuJvkbkDwcgRVgF5
JdotMOF57XUuRxn0CnwflCmppNJ+avzj+QESSPJj7Zh20KM6RODSJlFvjGiLmCxN/YLiuaUSFROM
z2CIxKb63Cxo90KWvTT1JCDZzzwgpAMgAL2Gx6zhHaeewNIkMi0wwBlT796kU+4tAzUfqEaM/szg
HrqLeOhxhaD6Upx7kbTNcd+gZOBtLJW3CUBA73B79lSS/zEhX/xYyuDZDB2A0aRrqVmbJcBvFiG4
QZh27utXnj2i/ZNzMTLvo2D34Lrj6/wl6e6CrWZFV6xZCk09/eq6KZsM4vOqmQ6uHHZ1XspbPAnk
phbuDvRhGltf/FFbfUaUV8PwZ2ozWgblDilgLDTHgDdt9gugoeXGXoSzFBy+yi0QMEn+/iwwjrWF
oDXiHm95anJNRUOEZhhr1CUTdojJQd/Hw0E/5+CYZRoo3FTvXbrNXSDNzAULCT6UPDuDH7jhq/6z
zEOCOBKzDpIm78D2WKh4aGfPhwVwoZzIpbgl9eNRfO/tI/vjrRFUkjjCiN0C/h/73TtDfa7xCt/y
BIYYhTKAdTpz8fwbFmMhkKWcz54QP/KxIB8b+4O03e6Xk5Q1NMtFdr1Kw+eslyfCCyKtOZPI2Y/1
VhGn1/0PcSsWnhmm+2+3uIsiroxQ0Zl+PI9nXE9ZSIUxVMVTBWy+/TTbA2cQxO3N0DqUIpMZfaj7
dJ5hrmWJCSAV3f1wvgJMbxgpFFcRi7/Ev8nx8Rv//d7jXzjj7sOB0lANVM/wLJbwVeXeC90MRx57
e2TJ3XguF5zEtbkaRsYKI0kpsj6XkYWD6v+gnoSPO4KV4TeqafkaXA/Com0aQo54tgnGoT+JvLE3
+4tCAhS3YCatUkKtwz2hc7eTExuu7lAn4bdHS7+qAzT4vubDJf8UPaIdrAQcmlQLBZBNYM74o0U3
gEtc3MLyUKTwcKkPxUiq1oDrFIqPhI/fUTCfpA3etZ6+HgxvF+TgLikz9gfOl5IDKLg6wW7hlQJ9
Gd/tJ/jUapDL5D/y6hmL5dDMF/R6KngkFEfWvAr7iL9b7Z16uolXKalllzcl0XjIkKJfLq0S1iIB
wDo/4jtIfwgckgKHQo93s62A5/Q4LvrASPpMAjXshpMvhBaku7xDkqQV5Q/IHiVVtGtR5Xz6Z5he
9f9aaVBxGPfVkN+wOmTuUthZcYeBoLPluHpIHcaxNSfNG9X4CvLWhr1jFENNCVSOP7Wi9mH6C1sm
qK6Ye+k5jY6sCxRQ1fdQNH3LvRttBmgEjjSevDkUXvgtSq3OBIZuo+C44FYp/Sa17aRKfC55oSwK
8SHwrA8LAapzv30cscWxGqqUuoInXYpsfgBckrEJgrXeJEPcsFj2LeX1O3/6KsfpKfXbKhONiWiZ
eKjViu1t0O7GoHMj3dVLnhCiAKyx0tUI5r/+pt3RHipkMG3+YB1Bn9yMBwC07V00LDIgETgtt+hl
g7bQA234NiAGGkf78MoNHEMayfJRG73YGz5pbNp7U+efRFixRrnaHjT7uRR0SroLNjbduPwMQL7W
LgQ8nlleDwl44qiSD1lqkxSAMSGDXCSVGEUt3+Sntw91+oWOnEibHPsgeELQNjZuI5VGvzFi7naQ
vmJMlYuutRC9PuZkCyRZxY+CPKuRZ2OX9LfghgQ9XeHR59hVCb2nQbqR5nOPD2rXlXpzgKmI0YS5
NVulhe8M01I3JG15wnjqRo/6IrAExvxZHXa3LWNPIMX9YioOPHT9L4Z9JB3sM9qpu34ysvdIuFnX
HvIfvAk1TIdWjgUlZp4lHT+HTxuC2r0xv2Tha4hZqnbwEu6DPEcYSfVztUI8drXHXesB5OKdDqXU
2WDCgMNNdJbqId4AN4XiN/MZFS1JCgcrm0ejha+vXq69NIR8Lo8EqcKrMWmTbQyKZGw5loQ1FsWS
xA6UCwzVgW7Lo7vwuxYrG9wvrIsWdfdZmfaz6IhJm6kXowpkYMlDIFvT5TBZJLOOAsnpI2rv85m6
hWTT6H9+jFNoHAQOsMQV15UGmvDlZEfApjtZRTqMfHTot2oxl73CeZvDX/KFKH10jtovkZ6Bd7Bm
92EvrPCEplRBnc+kaua0RmkSAmc0u66EtpPimJhEM1EFHALEaTIpYAPjGD4+vsAuM0BUgFesn/mU
X6uJbvXqSzVxo+sYKTUFm7GJTT8TZpWEN2T8aqr4SiPndO528KVsgGT6lwBKWTsWhs0Jana4mrmX
Mp6znSPlcOg/DgMGTuGT9+ZGxQ9j1myeCwOQ90RZim7+loYFZ5676KGeY0As3hmh2l1BumYeIsKa
WUkqVKP0npQakijncSxwYep9fcAXkhOqDoQyDOgOlghsz0gjzgtdbxQGz/jbu1ywLHwdjg1c7CIh
0jWb56WhhictSf+SEzuATPl4jwRcBgANolwVNNsf4RVHK0NhIEdKxSxKrC2Km0ZT78B21Ehe+A/S
IPPyAViOyIbz6Zphber0q+5OKPcbgUbFAQzkcGXNTA4oVoK/gdcE4l0A4F2pzhPEhYa53c6VOsqR
wjaHEKs0383FmAsUneYygAZSDDM9X1gINfPj3bEzS/4dwiYSqT2wX+lFvVgh0FgCIh1WHEoraS+O
JLH0fCdl184GDDIzuyD5h/T8wNddcZVOTklRkaHADeJZxql4e2C5k30fiulwgpLn0zQBLjfuH99Z
9ukYu7834uBV491xiQWLRCyOQ7sFEfzzl5dOtNAKGgCOCPQ2TJFQ8s8FDm/sU2CnqyOCnV48jM5X
tSawl22RWbQup1AN7c/5f/rkMB/yGIc2EH4j/JYv2Fxt9Pubt7a6HOTzgXCCYRnz5j8ED96SAMMP
VQcinZHgmlu8dY4kVx4jvcLWoR2777cDDSoiqHwCmhhd6aL5oJ20zbpiHxAVDnYNnOt7WmgyqBsH
ce8vrVfrQkWgj/o6LmSQ5vzMj9VV34leTDy6wdH2klpnWDs/oeJYegW2jOmDzXPk+cNLWf2uHN4a
kB3Ee0thhvHaVRImwaseR3O2Lb82Q08XQRey8YTZmiyuCAKadHEyVxD3JjRwYzezWtBoMbqS1Ob0
uHUXndV/V+0x2gbzVsjLcDwi/LyK+uejls8i756uwC03Bpt+NFrcd2zOEhQMEW7kR0OZ+IJ3ATZX
mW4t6+S8uhRyfqJ+OnpX36pwpTdUUWR1cq6tvcc9EW62MR3i0+IJXRRRqg6XkObkbTibXGOdWexu
Nl9OsiGTM22JAt2AlkeQ4wKGlZPerHZmfDa7nvDztOQCn5jIfUZG9KTJplVt0CDxg5zph0GmbOdk
hYKT824U5jo7pM+thz1875TUW6hltnKEyAOuAOAWCcvv62wKPXh+1BFMbSuyopeVvwzzbaP2CmiH
xPAqK39Yeg1KriOlS5uAfjvDNin1R1N+3+XTj7LOV+Muvns92V6QXSFGAlDQ4/e2Lvp4Ajhf3NJD
FdUb66WZHiWfpT7XYlrHPOnMSuy4APOTlOiSD3loBEpsOC8clj72CjMFIiibZmz1SeWOXOYAACKg
pGw7Pi8QNDhfE58LhqaHk4RSB1ykSeGgJH8N6oQvmRw9a2BA0WjaYhEd4zWkgkOqfNroGW8lkQZs
01Q9ulNfSNL/+kHC1VmxB0L/5ELS6MiWm7W1nCixNabIBe5cd3Or6YNAT/npre+6NUMw5hRpUtBY
VaZJDwTy6cLKXQRbMcM4YsCSHsVejpGRSu7Xq1djUGCrZZyyfAG+abqXDjCkVL+pboaxpaufNlCM
APcYIoNRe3118eVbYnMYosj6pm8LJMghB8jqvEbqhJec5CXpJAyc78QkrF1FLoyi883Zw6NoYsLX
KwBgQRcQH/bVbM9+2IYQlFEdt790i5nKYaoCpfWOTgBJiIh2Q/9w2MqWCNJFXxQ+/Txuj/qiQSwb
DZ6G6K4pB09s1tZ+EdW65c74pPBNA2k1WTRmKq05f4+Gs/WWQgrj5poN7qsdokVhL/NGrk2mPRwg
t8AjxkF+m3skIkMv8X0M5CC9y/L+eEZn2DQD0ITlCtFa8be0z9F/80fLWdgRzS2gpZGU4TZw5q53
jmRBhZbWFz+fQkEFH8QObi47cqY3Ed3os9P+ZH7t/KTFJbmwW+VGmUY+jzmR7ZBx85ta/3q1+K4e
K7yAhz1LNatZqdqw7Y9kU6QK+CAb/nzlpZ01sG0sIcnHfMIACsWnphhigC9NKNUO2dRGzOuuKjdE
kF80o99aNUvHSy1mbBO05PBEfH22coXRLw45BPGkELVU6rVPoZAv3Ze8mwP7ZpMlZAYFvbuBHFRh
pbIZOiwCHnjgjWRxqXqeGq2vfD61F0R4FtqJY0aG9jcq1uf/WisfwjAKoI6ktkLsCVftvcZl7Be9
Hc0cqm3JjWy1T8B3r97IcOrrr8cX9x/vhxdaXEGnhbiLzL83PaNXcQBGH3wTrb+Qwgi2PPPrAO0a
ee6OMbY8KaRkjpEDB4YBeyQ2sXpKtJa40fmLN49HBn19nrHoSB7/1LrrpYBzt/6D1abWj6g+5X9e
T9oRpVc7cZcbo2VjLlxPoe/vKvm4f+sae+IW1XQxWik5G5HaWC0MlnuUyl9vLlkqFuLvXhZksuuu
HtIZAIs4+zrWj6XNRzI+4cXmtylIvpd2CprETrJ6294fxt7lZSVQJkUJ6C2IIpL1UJgszt4Y7+Y2
B2e1C8/T9GdAl+KJZ5lmQjBvL5N34TRtRj+08YQiTCjZOWproqToxK1NgB99eAeufaEGbR+PCx1W
1a90OSqYqOliRZrMXyQ4zUr1htJZar3xYT92deJcAVbmjwYfFdNKVx3zRfedGbaciBBwG0tgYJDN
haWa4tiKHIuHGyYfCPA9+j1nlM1L6MtDT6ZmM9r5fWRKZmVZ3xqDQJGPu0eDajdxvfAa64Kjtegr
4frbEXjNxRLf9eUE3LeDsocFXMG6pz8Y6bg+K0YF7w6rsB5mhkCoNHO7LwrQHCtWt5bOv3g6VJEU
8/7+iPhWxARp2StEybFy4dHoBeQy+wf/9OQKGr+UzzC3BRVe3rClCAxRQLPg+dD2A1DGTD3WPv+M
L5QbaxVr7Qw6G3FTYW2dnC0taAQRkTxFnvzAyHALTVin6o+xlZg10xNFuK52hdN7YebXNGbulPC5
C4sVSpqC3/rAjTgF66BJKnPIN+ecTDa/jqomy2jFWNPVLpxfIj62F0C2JxmR0pHqWqk2tgSA2X6o
/hvh46IZmzShClsNb3qdbfx+/HSaSVNhAS5mg5XimiWYbMU7AujnlVmZtOvt6nYH45D3xtM61gLV
fAOygPqM+6g18IZ8o26EDls2XZmsLJwQwWBn1DK3+pf0kppFw3y+qtfwdfK/CIISzerD30KONrOt
OopoxMoB3Il1cN/VMm5qQaDCnivhgNfI7BjdGHK2s2nAbUgWhjzsVf/HOS5zez9dWQLB3XUyZCFp
z9pi33XalRdVS5ir46PUXcSOqTq0/z6uoRxx6/qX6eC/5xwFux9NAR7z9Oc/Ur8dNhYOd0k0FdIG
uAMPpaXQfM0d48XOK+nhY8wYRjceoik5NRN6Y4bCV9fHY+Kb136C4LXdhHwWryI3M6Mz5dvq/0vs
mvMk6h8BdVgRn1KK7NdMSNHeSWV2J33lU2gv4ocUoG7MvjKloS5UMf58bYXJbhrayUvh+Y7i5iVN
YZxnLae3D1iya+lMd9EsLxG5lvGo5KDvOI6s825s+vdyGnJJjKfZc6TMqSli5ugsrqvj260Lrtlv
oGhRmD1FMCHiVJS7Kcou7hoPi59VOzZSVF51u5AGfKVdhMAI027yawR1d+aVc8EjR0ziepdWgtiU
PMSHOWUb39AdZqCKvEyt5c06bXLkBjnKQq/aVI8FjB8ey47evUrXpA5IB13BcnnswcxFuA1v59g7
3cUAGHT8EXirubrMF295vAnoBQwWeepFxplGNBqUaczvoGFZywoo0gadYt4kBurYQHbwGxnEfV6/
YmjlDgG1CXfLT5odFfAsqo8hgNqd4qhWKqslSbVyrbudWiRlOinTIHNqg9Zdiz0PqSTGRvJuKN6n
TLtIb7s47wIbY4V1xNoE1ZfuMPUHC5MBjdSLV2OmIZg7Nbd+UOmyDUfC0Otme4qPbRI6HS+Rpwpc
hK383RliCPyNEYGCBTGV1gvJIrh1sjeqyM4vMrutwU8+HVpNI35plxlOHspVJW1XrbmrS1ww6E5j
5BLLY6MJrN0+unoNLnpUUfKZlxd3XAvyU6VfWuanhPuK4dFNK9YGBMwYwhsgoQnu7aFfSCSrGU0A
QdbJg8MnM3/2yT4yvTC0L6f5+nN8FAUss5RbX0hvNP1BBYPsLpQ+2H/3cbLeFLOwVHvpFEixbWG3
wBd3cTlCiHZySUHPGrJtwyJ2N1k2SCRhYOJKhVpFNa5VWXmj2Id7Dk4aFCGIJo/1sEuWJT3J6uOJ
PJSXor99SoadgpQHbCqlZgI+pu43NYwwutyphGVdXLcELIdFfn93E3gUUtsKeNhMbIbBawHiEVs7
SXUS0kkI3foX1r7s/QcAfD3F2yfL7ZSM5qupsKqtBXk6p8qeSpxTh+5646B+r9mjK5jFW9TGRPvU
iJx8yttw0+1j9WaVYr7J2WpXeWxU+CX2OzkMIpgrrasTGtduwAbkjcVHe5amtQiHPb0XbG8YMr5L
IZsfK1gBXxEv3zQOibARJ7Qge2iK9wekrIwKZYsyZox+1gSg5LhZhC8LaWrPOdb7zur/PLZT9rCK
5z4asj97X/znw1GZbBJ4xJZ8XoBsqTJLZlUA9D0wZGwZM1l270M598jJCQ6avZbqdFppKpzG7Juc
OvKNa1g37M2eidgs8F50XuOMyfCd1Y5gEPbZcmUXTCv+pZ+B8c6zNgCpZcXxHgKqC5vIWTx08mPK
5VXFDmCxo68YHGJmiiWegtTSebKQHADmaa+xtvLdAACeZTV9BG2kqyu2e9fNtBXz/2IBbYCTCSX9
cGD5OZIXuGD5fjdgauq/9lSVCjuq1F78OAnLvAtppO97MZJdO4dA2kaT+7BVcHSkUacLFITxp04F
IVXpWlvZ8Yvpx/BwMQzVC78ia1sf+ULaSPviumRGvwSPM2xsEAuaQxNDtlxKN4XOmx4t9rlbatTK
Eo3wBPe7ZWWte0DzEqMVQ56OlV86lVI6q0OGZGOnIgocvXNuNEvJjdLc9K0WJZ+2Yz4+ky1moZe8
5Zzm6yJkiLRpYd0Vi9odRAHs9MAGFp2lXw6XLzUa/D5dqiQqzfRb7CHpr6vbhqhlAB10WByxG9jx
gRKf5+Qa/Erd1LMJXQXeDMn9mJNGS1QQGoHSC0g59Pq2ublBwRwi5FWKvuf9ChChHVnyieyhLmXa
74QBYK6XP6/Mzq4us74WUm7/84HybbOEhLLb8a2DPY920jWhjizxjOK2n4U/GyMvT3jKv4YWQQWm
+jF9P2xRjnadJEg+q+CI4iLQS6XfF7LjVxlyvL1uGVeSylAMySokNBX2AWG4old/iE1NHxomupw5
OaKEYPHfN5rAc5kABbJG8NIpzw1dWWNbTucluEonq9Vt6VwJAmF97wkhYQXUI3ocjJlyRln1tygL
0NBNktDdadphfl6ytLOc1SM+owyFmtlVzHv+lVVJ6JlWmaUYI2VWSFu9V7/IC6D3rB/Onk4GLE5X
pEhb14LBqc1U+jBqxIs7qVGN5ljnVFzE9YEvfg5RSbnjJ5ujqazNfcCCjc08rqK5+qDeVwtgYmcM
QBP6WkRe3XxK7XADZEQmQoH/jMozp/6nTf0cVzktytCCl37MT4A7V4XqpWUHVYUxL1O5twSVLdeH
r9KmkN3WhWcd6yVB56rIS1KbzEhqnlgIgf1EoUcYQcRyxTjVCyeQVKYIyPZtYveOCqV3oIO/Jv8m
eTialDRHz6GGii43pMAN0AlGEXgovd4LRT9L2v7L16g8032ZTRDabW02bbHmUK2augtpAv1z9Iwr
dTigpQWajjfGvEFJonkQeeE1pNNr0qRagNT5+zxzdER88KSzA/jL5GWgLOwzsDsh5UuOtC5OoXjW
17NwO1j7xy+F3GI0Zqf7UmrMzqw2kHiayFwVGebEyEfBkU3ozWpAPcS9VnnBKKoBFAiY9bJK9q62
PHwAEbro5ELbJ8MUy3EaRsqvh2Tb0IBFOHWb3vQZ7X0haQS57sK6TFFSS8mMbIKEnm9/xXoPPs5Y
8HfOdreg32DVpwcz/Oq3S9ZVxNeYGtOD3PLNzuIyz86wIvDjNC+2tLliufviHYgKL9cOqA0qULjS
f6mmVaD1fFqH66DmZ30BV8GWvHYYjwQZENu2R8PFGa4HK5n4HKtyxLjq2A6gAlki/vW7th4hLOA7
lKh2RYzFzUs7MMifJPcSrjqs3MP4WoLFdcI6WbSqNMqQQ0NOMH7yIlmP04br2UO4VREX00MEUC9V
2WigPKe47x81cOMOsnWE12WGgfI/0OCTI0D2E+YgQf6NJidyRNvI3ZPT6vAgg00n6/cHTEkJ9xJV
WTLkSb7GkYWZt670z99g7JHYI3KfHHsZ1PvHUm9Cy+qQrDttAy+JJKJbBjJXqT5olKIGUnkHbppD
fe4bWerwQ8d8qBlZaIBQk5prxh/VADYZUA7YpzmiJJ4M64MeGn/tM42OcDx7i6SBg4YJ5WnJofv0
fsq6qA7HWlZxGes7ow92WZ0so+XczRb/3s+84XXw82J5Y8KhEbQJrYkGUEnRGlJf3nUqqG1WD1ir
i1i1RaBHh/th+LkuP+/+OrWdgBtkGDuwOhnFPP4CdfFg1p6BnzhNu5fTxzvPLNbYLFZs11BFSbeO
kjVyqTBIfWQaIj+nW5eQ2eceIy4SZ8U1W/sVX15oFwYvdXDoJNiVI9L1PF7tNshrCS5qft/NgB4M
z//H+hiPdkD+qSXVecq6vhsgKlOY5QYTkbMgNVxFcMyvaMp3YO4iVBJSQzXYFBdbd7NbjOHYhcpL
Prz5rMcchgopiF2jQCu+a9usNqY2cZgR9q7P9reFTaYlbNg3onzGxdXWVTcGDOwnCPJczrk4hs7P
A/VqmNpvOX+ZO1IhX7JfresXm22EWVGPRO+gdtyPHjjk4atYxqDJhsytiHyM6c+w1GD3Wh27w/qO
GHQeJVPxEarbRIMVJfGzGH4L8Whpi7Z6tiP5YjwPEX4DORj4DYdTSJ8jX+ukO4F+XwobYOc5dBS0
mjm51Dd5oczCVd9I4mmXbrZmur5Smm+8I1tDUUG3SWr97GP1U9RCAI8PS+SkIduUzNENg8sXPLoZ
efzCNb/b5lPdqAuQvhlBJPC1P46SdeybDRbdABUIr7hNCAdkJ3Rn5IpJgq4gvap5Ex1ZcHShWQmI
YrBI8BD4cYYqv6HR+Tuj9xlpCwJpRw9EMHLMLnw8ilL1V5hhoKvNA9NHlksfPpzX5pQOl4TVKJSR
jfiAsw+IP5aVzDrqayAmlTcSrQ2PD52d9UG3qJ8SQUr55lj3SrMK8hn/CGDD1kUwExzTeGgKZFZQ
g8VAGHUEbTe6oaU3Bxa1SJhWda6yOJwVb4CeW/aLVdwyCImIYf/0JQZ6FLQnV9alhFR6/Bst1eOW
hd2MYQCHvyFvi7njucDKNlLXWWx5ihTHa1e4e3xeXj2qOkyUJfL87LYd/eSzPP0kIrU6aFky24IH
vgjPTKoSxd3yFTpqjV/xYW+mlZe92KvGDvL+IbZ6LWC5H25bn5+xF31cgziwRzKyhTAwaKMjfvTa
euJ+H9q2NzfqD5Vdv2r9YHdR2A/k+oSzjpfU+liM3xWphO+uL38qxO7F4KT6eurwdaQs4tmeDelH
5aCSvwRy8UJaQVBahPh7jQ36aFsQOvfWQPr0nJPKQZW+MR+MdwfjyTWDYXtKjEjZrStqmHAKwrkY
gpxdYo6PAvwTEQMOyORJn5bU4OKV2W6hqDc38aCPElc+FYzYJI8cIEm6E5npZ7hAd3G+YmUyIQkw
nv33XnqIVinyzGUJ188Rfa11WsIx506IV1oMiXM2eG7wb0BFwbkUOAmC4ieuJCGCnUNbISQnpSvM
9vvTIvdKmqDd4d2+R6VY6kcWD7zXQUOqD08EP92WyKpjdnUfqluff96SfGAOj6vDSKkxf6cfOc+S
eGkIYU0B1HVKkfKajK1+HVWJu1We8QKGzHkk/GE6QrUwXJEBiYTsYUxZ0Lsjp2ZVjd/vUlur7Hdh
9UOVpSutT67jAZk2Ad6+UEUc2l87K7Sx73qNphn7ZpPK8lyWDmGTIsAPBVJMURKnccetJncxiJ5b
bWAEb0cc5A3h+F0reBHV7P5vhTv5SpvpcDFeJoL3rPQZh+ppUnMGXzF6i/1tthdLZ+036ngBzjHz
A7cGER7MOgPoA2VZucc2To4dy6VIV4bhmZlG02FCKlg2JPZbnAQUYoOzgpNnQ+VZk3iAvup3vXrH
1YBm+dL4oyaXUihN0h9+zgBLIR7xVsZu22NGat1VhMUo5KXfi/8Tzq8SKGdrEccX/oUL7A7VP33e
Mn4uPNBWL3EwHx1D4cV671XLc2V9TBXfDs1Wwl8hLxIzGgTpa7/XkZHZqG+vxGNJmq8xkJq/98no
VzxtILIfbF8E7PgqHvGg/jUu+0I8HLIWDLfvS2/WcSsbmSCppqzUb6rGmHPe79b07Mp2hXH3L0Fo
JqOMCbCT8EHaYcoSN/om3237QFDuO1iqoNOqlSAs90EQpuQ/BBFLc4zL4MEJPZIAUIJy4UrVkCHv
tdXR9IUDwjNc0hiHjwK6ZPbkFeaCm8vHqjp7S15IfyEoWQXkaBN7+UGmn+3zeqIiC3GnnnJBclGC
rtfoKpfMyXPIEeSmuzGE8qdHYNGodYmT7rweI+SzsXUvbVb/ykhqjLEDXvWow28jYxcYqyXmGn2g
TwaTF3y5yObhxBQ7COZFv8iWXpWLXZjK+5LapQQQWW9jvHeYNdeK4xAc7eKZOMPla6spJ7MmpLHd
Oo+M+/zLnkjK97YMuhVMjZ1yEp8VU0urEQHSx5yCsyZKlmZrKUHTj5534WQ7RXarNUBHiWT1G8YD
4qi5JYZVvxWnxC7Jpe/dRcc4lxjcGg1psE+PFQIxLQXNVtn+B3zhwSUkkyD0TTy5wqJhBrvManqK
o/O88MalEG1Tcu2uHxPxI0Nu1ackHgSE1tmodwAzLSGbSkNN+irJlPQ9zpL4YIvrB3kkZr7z+Kop
nuGNBv6dzL6mBXIvVapnm97dnHYCGaNcwZfusBLqgvfV4nRcXEwvRWaowtpWB4lNAMMGjFpmG2OC
vCYfXEBKXOmYU24rKBr8CF9BYwa9/SV25aKNK38XCZuRlE8I6J8AnDJgEej/6wA47BxDAnHu0cSj
Vuel/i3RYa/QhT3etFe43WoWyIUxAoBCO8f22LoiQezGeULKDh7sz2aL1edtTJ5N8+G2dueDR4rQ
V5dRBKSiMp/7a2p4mES5zfDpjgpv/+wV0dWD7KKSyfOhggPA/S+FCXS3ylAvnrkWMEh4JQIGV2nb
bhBpVruJlYsJFOIoXIjkIV/3A5IcPnYLEmkcJqnR/WFK+Efb2/mNwZTWoZ+fY24BwNFl54Bph5vL
42MTZhurHjWvEn5WC6c4vVF6z1PhcQmFox9zCNw55lYW+ZmL2L20OfY4alI4a9tEUVQZWlZsvkuv
i4qhZAcp7ynFBKh10BjOx3/SvwelXnxfLEabUVwOdu/GpBv0R5R+ss8fWYe9VsdI5uFApy0QaC+y
DI1ZpQr+LMoXkDlcazZfHmiY8YKdDOYgCQE+O8C2OQ4nLx0JGHSN06y1T8fAeNgcr6eEnd6tY/RK
NqkUjKyQ+Bz7PaHJueO9IEzgBDit54+9t03qNEDm+s0/HFi6MvdfCBz6yJRAzxyqdCNwrz+Stw1o
MVaGGjPV++r3g47icMRBFFml+/6DwsOnkkobq2vlGo0l0VtBPIvoOjuT4I5bvO4vjE+yqyFnkykY
mkiZY9vfT1CWjNRYXLatI3kH8TcLBxUxS0KXB+5/0BjAjWwbTyRUbK/sGrjR2h8k2hyGkifgMTL6
t1vwT0zfEvGEFNzAgc/ZaeZudbuluCXu/Y7saQxDZ7IOCbxbwBLF8sX83TL9iJsc3vLPYU+Q2kjD
+Qyrs9StzZRXI4n1zTS6bzdWxvTHBqmALkw154xEpd06SQCal/z9TwRZ6fISDuSkoF6jn6wJiI05
OOx+dmBfJTYY05aC5IjVcm0nCbh/UK+2a9FEu8Bk7subDI6CiFb6aE6p5F53GGKdeXK/5YPNtkpO
9/sU/devokT6LW5Vo0a2IFSTUG+aH5hX35XHUaEW6f1+NkLe4UGjT7mYrchI2vhnbcX3Qd1V/pnr
kWWj/AX4YIGPOlZ+yBn4G+nhtGKAuCVfsxjS6hjsDEGN8LiRKrRhu2n0TZAgso3Hm4Av9/W4fYaT
Oh/bhFW1lNuWvN/H7LnJRBH283Am/fbeapepHwOZWroR+wy/QqpjpfJqkdwdv0GT/hJIUJ1RtUA5
dozG0uN4yR476rF+EFNF3dv0FOpJZ9ZX00XozpKUr5DgBTEaLkXh2+sm58d94m/gIZ+0Zovcb740
rKrjxALk6+JSrV2PAoPO4oExiLN0mvhaZLdZuX3avF0GU9dSdwrVGyVSB4ZNsIusVGdyocowiJcZ
CkxcucQDbnp5e4tSXh9GQxsrFHxplifNz9pe1DxONbpPF4J0sTPj+ulYAyx8MOgLAelbnvZYN5Gt
bX3vxRFXr81JmljP5pXA6Oudr5m/67L1uj3VS5RXW6mwO46bmjM/C/4Tr1SmWoSYUZAXLdb0b0E8
XTi5SlTDjG39CSwDW3McMJt7eMdgPhC4aqcThCbvSwo4Hj902S5U+6cGTZ5WR1vCwEox/yKOhR3J
ep5ad3pBauULfXsQWzKptiu2TXc5slBe5gC+BJBGbmx172xMmWxUYh0KS/FOvChIFLomWwHhwPCR
F9shN8hs4E7L6vuWz691icBv1ZPDpAqJhZ/luM/cSQMWf/WoaqXOWWjMr++eUeoPkBXxRGVmXgAN
VMGml35reY4OzizqZf6pz2aKuWqUzpkK5qTHc4ZziwM/yej6MMETO4m4sJaViy8cs7G/Ca3chmUs
3mb4qiEqVEaDC5OSf6eqlcDupPDkdm1aJ42Sjktok3YhARvJaDh4MmynZACoXspcFbp2KlKeCfdZ
+3Cn45GrwK7XkSGvU3xYiruU+tvbQJbaoFfZOBCJFvVQz6qxplalp2oHXX2ikHRyZvXtaOZ8USj4
WLSxf5Ui0C5aMfySorV09cKYkcsrFLlon3Isj3DJwF6fZCrWhK/2d669JZx1sIap2aZGyeCv5qJC
dGR7A/Dc7JVgGlN4Sq6d47CU9Q/S6ejzMbpYbQVdWyjV0FvTUZzEZcvRdIaFTsNffiJrgWTDsAmL
nphop0a/c0mCHStCrVoadn8avPW9e6FnQkBPf43LXkCTc0sjvOBLKHYCRGVDiEbf2fIXYpTsvbXm
pZ5gaqlKKV+BnDJ5bECtMmOalcHJk71GbggnLEDh8cIeNlVhDkqJMQ/EP7Q5eoJQZZ+ly6l2wi0T
nc3nM6a9K808bf20++Z5q47eKSFGAtrQRbipSZImaAXzL7zcoVUrIwYNxqov3MILhAif04UUltwc
dGyRTail7x2GY1EqNx3RHSRUvzuy+3IKBtETPK5koz81eNfeQKmjkYxpyxKJJvdTDHaGsIE6m6uk
zzofiWeVXNiKrt8dbjqtMf9Q9oH0WAgt4CzHD/VHi88yKJwDy3dv0YdXZFbp6bwCL8LybbYriKkW
8LqdQUUVqsLXpug7zXBkT5m1bIAI/9ipThjpMevYPxlRPWUPdwvuXDE6FGyuiq3p4fMMwxkzVB7M
DL0l+26IrPcVNpVyVdiIJjWEmfOXZPys6T5sNVdub3OxGvr3Xuy3RBw0BQNpeLNGAaWvY5G4hkca
GUiA8kgOo4bdm/OgIOz5xEQUhL6QptVr93WPrrW9QLXTdr5v8sTo14PPly1FME+JVE9ZVgtu6HJG
rDQ/2xxfm0bWDcfDJYWPNDYrPSoUtTAWpFbELXetl+TI2WWvPvj6ijkdXwusEfHoSDeOVel8B5NF
GssqjaT2W7kkQ+KA0PZ7nVZ26bMaCF8v/Ij3g5MX7RH2iVYHMoc3rvNXikmtm/Cn4dTeaJXB749S
K/D2Sit9T8pop5jZmG6hj//u+f0hgihy3VlOH6UleI4SQOnSwq4C3e2qmJCRKMEVsahUr0GDF1Ek
0TkVup8L6hzKyc0jipwbzU/36F3uhKq92V6wYZwaaa0XoZxB7sLFPQPAR6qVrdqT9D40CSXlQBBA
gzgk0uJCxoTqL19b45uUqiIMq6tm5iLaEpjHTceHzzy44mMebVFJ9AO4DAYtq7QL0GumbTFeLz35
jbJjpUbCcBjMICOj9GhTxryQEm5yaN2fwPnVCYDvf+FwNvdp3hYpsLxCIRn7+y9IjuBb+NoSMHvo
a0+E/A4s1OhUB8ktYlZ19UQmmKQHoGE8vXJh5ITK6m8TGD9TtbSnQnliuYs3yp2TFHRpuKo/XXAF
qqcdQVSwJeb/yI+Rs4h78WehF9VjAd3UfHppfInO/Weh5EctRvn+CUR6HqUYxEBcIdYQ2u23ymxV
VWFbboAbRAKY4RaCLghLO4jUYxXPuRy9EMsXrT7cPFgUex6KHi91PQDWLrCyPnxPNscLp0eeJsx4
csTrTuqcd69B/UXI44Fv/iUct4MYuPmAyEX1z8KWkIxWGHKP72wrKNhWE8Oo/2i4dHVAXNV2FaOF
DTq6vy+7jubfeZBNJ+IAAtDEP+nXKY/ps+3PxUDzQvprUQBoxnZrfTRN5wuKtLV2r1Yk2Tj3fUqu
eHUrFGZFJryzPtImtEE/cFPcjpodXbnSr+oYPaxmGuzSGL8Eo/mwX7c4U8yNeTFVDY/dZMzF6Y0K
Yjh4mMB4p0VccXZbSKBRkMZqrokOZbLbXB865gkjucTRf7U/1Raefpk3kv0mA+jp0bB8HjYi0Zyt
GDBNQAt24SG1BuyG3JuZD/y8gvNRBZ7t8VjfrNjAklYSBNAqG2wEupCrxAsqWJ3TObSaZpSRjFn+
HXMKQAXUTR9/N5oBgvaAyLjFLzu81tiAq+JgyQHjbhm5oXfOVKzxawll81IdiyaEiBR3XxHZHsFN
COjpAzSwDtEG9oLyEHLBVs/04ToG6gY5K3YggqDUn9f7AN3wTZ4j3sAARun+5yIB6O8Wrh+klqN8
nVaE7VdFtGRumi03yyAKmLrxP6ogKwdt4BOtudRrg3MiaF0IWS+zFbmfrTSc6BhK7q6RYBAduDWj
lqEvBySyP9eGu/HzHgA8FYiVYcRMghkiI+az0EW51CncrHs7WDOowWTatI37++LMmsx2UiH6QwJU
zX+1FTZ3Ak4SJB2g+m7JVg2t2wD+6R2JwdmyfbOJh3MeC11hVG6kbepMjzF+Zuj2hVnTWWd+aAEg
FO/BjTc1S5TM/LyVAiIAiNy6hUFOmNjd50rNMNx9IS30lo35peGIdNlJbf7VNUgcUEkFuHzlE1Pg
hiiJFaLTGFcqokLXwEfez6tc9iXwerI/Ml90qhScfABus6maNuRX72jeCiTNOKJ1M0v9Oy4QT8jy
RBk6ikHetPsfQoz5BO+iGS/6b7bTOqjEKNK5NFHLCRpXgoQbACCegj8SXHkuOY+uDsa5SZ5BjFb9
+SLc2/I1vE9IzQ7mnLTmOgnMo89k4kds83DBby0BmuFQbjVtUTWC/BG8hPr9FxSLQZreGhHg/JCW
tVLFnoaFOZMz/YJqbjXeKxWL7boIv/iI+p1p14KNOweqkQjDLUyKf8LGGcboFQDzK3nD4bYJJnSQ
IWmfa95xQLryUkwDmiaClgBYzs27fZSt8jvCSxYFWjTYlMS2glDkIhW4QEGg36SXg0KXElNYF2Pt
jScQRV83jMSdxMuOoWUur5YS5LzrdaujpH4m19FC+Xjo1CcnHUfjnsYLb86gqSIlhaHabNx6dap/
4VbSoAXYoO35LCyoCUTEZZzX/ayfnXzqDc9fXrFWLHSC0FfSDaz/+FawFDYY551p9QBywV42wmaf
zZQCZdKejlcKujrhkOKEiEU0F/saho7gknc/lFn1axLnyysORMukqPRFD4WzteAnSupJuukXxSJi
Kdi86N7tMBGMfghC7obc/WcYlrJZD1PCVPxZRU9JfUCe9BtVI5ghZ7Fea9424hzmlmMp2ymtFTW+
sW6FFJS23dQG8SKrRQQn2DiK7yY9/mPWEHh/67yPDJtb0Kq73SfyKdvFcRd71JKxYGEZ5IskFLKT
QV+elJpD2XSKcN0RXmdR0OH6i9A6+rlG7Dv/Z/me/XSXdulUjotzliL2FZI0HmLbCEOFdkm2FK+J
W+TPEoYirLBwWGN3B/KM/4lo28bbjqj328dMyFtbYvrDmrZZe84IU0b1qy7OgBAJ8cFaOyKxb9gm
U7perBF9271xwEgG0S0d9GOaU7XC8pu6wkyOsKP2HIUtbusVdvVrgrEvUFb+ZvO6admAhL42Ea8C
nQ27yygSB4Tkh33QfmcHSpB+kU6ZW9nIJVVr/6l41HaDPdogOkvBOh4/JhUlqdefwtEDms17/80K
UYviZpSqrsk+GUdOURucBM9QblUPy6UbaejeIRoL0jgHWzeErQe0sEYwFMLBVNXGDGMTl/w0nAbB
tjrcHf2Q+adzmr2lclpcpFBQaumOOZQWLvzjz+5hZ3KyS1WjPOSPT/ZEvWX1I2WT/FiD259IizLz
rwbIwu8YhKxWOLXgmZevNwUq/woK/iSPL3AU9yrnl0QvUVHY3n4ZBlQas3pPQk0vef8yf5lHRW/1
WOPe4hd+xYcddzw6uuWU5Yyd94ISOk4gHLXoNoOsVBWGxDk/x/D9JcR+tzCmZ51bWvAG8ZWFSXCa
nFC9pjtdWTRXMQIkitpW+MEGiGA3FWmQcgvQprf0Tek+T2HukScrrRTbI6kZNcEF+A3DMzI+WTRN
oxzZjqANmlwQZuXpTk2aafXax9JLWL79rZjUgEyt0ZNh+N9N6kw55gyyN1vbNrFQrQLZdovRUHAP
ukHSkIe2F9rJSM/VGkO7mGNLZlkBk/d9jKmMVCZyt2DmehYxNUDHQ/InEGbaOXtQrN1SxjF/jtSg
JnLwzIUqw3AligZ4H3PdpkhBHEtxwS95ZspLi6I2ZQnv1lW32o5xOWhcxq6pgbXbfZgyikfu+Wie
ObMahbQgnSXL3phOCe3pwvKr+P/iXDjDvobPIt+mLEa2yEdoI/M/65viQ2bwKzjJWjkkH+yt0Zr6
SQpL2JO7Bkfp+XXyD10YMv0qhpuWXMovF9q/+Xja63RrrzHkB434lGdrXM0GvJBO3kqVCuOFkMnr
xYMVOrhqU116c3gJTQsqoEwD78Rj/6mQlF3D2UOOwtMrnsZVo8GrtZ6dz+qm0FH4A0mlgjm9t9GW
H8udftwINeaX6MciXth3h15FgLrlCvlS/4JrdoIq/Wk0ilf9BtZL4bPW96qyXq6G6i+pBPiHS0TD
6VUZMwM63Y0Tn69+VpvMt5rt1Rq20NXNMDdnbgppJ5cKpJZDtPTIkWyoXszxSyZFdYVWGM8LtzwH
NFkEN4O6rLY035hiDPwEBEeAkv5um1VmJjsiY4YRk8dGDvkEa5PRwDnVGnSbYtBCDzQJ7dSdAVya
+FWIVgWmomxC3orWYn5lP6jX280fQziBIdZWz2uYyYgxteEo/dHkBCOivPCIo1zJOeRwmWgMqJa9
85nYX4+WK76hEcW1Xol0yJG/vhptRXukmZlpJ7K4xQeqNuCxHbcKH/ckmlkDF9CEQuZGbdrbBuTC
YhwSAkKaLHF6fK7lHkSt6Ngi8qgtHDT3wmY03ojRl2Ske95eECz/lA8rqigv08ec1Da5mxJoXV3v
bL43OER+XAR059Plj7Qd3ixmwJOSmUuzVP2hY9PieLEuWwikS63Z8cLntn/+x5bXJVnRMDNibWi9
fADV1RouHYBYWc4K4Abg/I9ZQu9h5Qh/6LYa0hVGk2f3IYRun9KZqcYitlIVAEMRwFndScHFHCc8
WiC+QwiGlpjs6KNy+XlOj/OTWoB0g7ShZ/fpmpxBVYr56G/RYPkTsq4C6VJbZ9oZxrC5UFtTtue8
TGUyoNJDHL9Pzc/Q1i+TYKS3hDkUrbx+2nVAQcbYl0GuRo2tC2dwkFSElyMzFiUtWu/3HeL6kHQy
rzFENy1eh1ATRfDUihfqkrGSMq8EILJXceptG24vqgxxN2vXV2ruzw4R+9HcM9KTHBEFj6mh4dbE
S+KmwpvzTN0F/2/qKHZCL+1ZrUxJd/FX3pTr4up0LowKGsS3pXAaajA3LqnHxQqJIkDubuNSbx5i
B8uGkjTkDevJ/HK+EY4QR0G/1wAIXXvv6uQGSVxLgKYrppZDR5gmhFdGrCOj9auRtho3GHpjpWSL
x6r+dHDxtreq2s6zPD3FYfjK80/OMzLnole8h9phPU97X9poxRBDCYYFeIgSuJmzyLqOj/dSWWYE
uu0lxxq79r+MdZDB1w6CWmvllDqQIvW/jtrZHGn9uhGmywjstcnV5wqP9EM85oVRx7cIqEaDZKoq
nZ2L6+7nqZPXV1Y+t5TI2uiPp2vDsgSioxRXG/pgcmxELBbKEx3FDK/yJMsykQSgYVYzXrBb21Ke
SXlZfsQ+XkrTzdgxJESiYi+0ihImUQZNDhVoXS9xHg+/Su8ns9CgEEV9mlUmqINOHMz1J+JLuUrN
X96ESVcI4GJWQXxyeToPRk/u15xzO5srwmpyjrIJ4NfkPhvz3N8PKkU4ci+/5v17UOXH8bNCX7Vv
CCYXYIvtQ/dXuReUNrg0RQJo6f6t0hew2PqDWepMPR6cUokY58/+tJPuBh2eaxEdxMbORu+BJveb
Sc4vvHacLTkHG9DfhD4nfW8J5VHd4M3nj/5tLpoaarmctUwIu5iGySp4rAt6QmFLSBH71l8/VYG5
FwWqdAKkMAFujn37HXgzy8+MzWllxbuVlXzje1RU6kdi9EEfFZZg5b4m5H/knUKYHiKsX6i9Ss9I
uyHW2gdNyc1JjlwaCl5OMkjYiXLV8JxdWNexo5v8tTLdKp0hvIXQkn2FCGdsfFN3BTKUkmUXVDBQ
0Q3uPFcmOpXtUKKOzCBtvHbkf3TVgKSTHrEIfgMCNRCpQuggguPR3YU7qjFzJt2cq6JoumfMeafK
5vUuTgaX8zmkr2ca/cAo19KRiM6/DIYKZMw5x1oV9O3I3IQE1Isn6LpR1PGbA53MgK8+9Gxan10t
yJb6m9QmZdchqmgT3IczwzqIw2lVr/M7AScUEcVJ/jhC+D1OqmB27s7jcLKj6p/CjVF7GG0wABRi
d6e81bLMmtQ+/y2UzayMT/6myqXki1ZIPLZfgYGAnLcvZjspRTCU1idDNkoq0FQtsI8VQ+4UhPKt
h/dAB5W3yz+4oMPUQNEjauLj2MYHBUjrzhMUtjwRb0vVAi2bodB/vf+SO7BsGIaYrm/8F+0OmLk3
ZUKMayny3E1DniXuJ/7LAFpvk/nLTINWk022deXcTsBge0ehqWQSAEOVfUwYeGVtU1Xv+6FDqo53
2J2rJjK4vvV4EV2tAdm7OJvi8VikjrrFdmrgH031E9aPkj7P6hfX0CnBz9iQVjhssyPM8C0D+yET
92DyAApTnnEbqLbrKdbmuZq2A/fVo67B7PuUR8fq5LS0SPUFtWAaEcgXh9b/Tjr568AkLMIc/4ib
zW8uWnu2zEmWy2kp+t6hFsoVamPARTiy1hVbXqbIpyI9fKEWHbffv5FEnLFYsC+maFpaTMni2AhI
GiVXq5hwnQZ8BsSXqaBPBncSJQw91OS5/WaJN/hSsquUh2dHiW6wQs0dqCJUjASu5iFhyI4hgt9C
26Hx8Gx74EarZe+nhUQU3T/dAoRepwTGSJzKlheHHMC3+RyVpD8lmH8ECNx/Mx1opvnTrjDNe9Ql
Qai1UKiHhM380kwrH2jRqz+0JHP3A6ecmDmR+Ugz2ZF7Rj8Tmz9qCgngp8ZAtLuPi25I5LWYKzkJ
Cjq1JmJyD2VCQ8j1AJ6iGWe7Xo1p0g8k7SM2w7kOlyh0NcjzXB15iGgBWRD1XEMAKRYixzwPrZwB
ht3QCAYzngFrAx6cwMMAmG3+Wa4FFmBnjI4uADPW+80liLBSAifQSFNEwgVXWDZALO4oq2dxXy1S
e9RljySXRCmdNCkX/Xo2N67Pl7e67alL730ye8FuK53XO+gduASb9LvpWyx4UXX/+YYex2UeD446
RrIjhHittk1MeUhG8hlf5/TjxhnNEIUXQJ1FgMKE6Qdr7lxdb75ddycxg7stC+o3TMlPrFuCViIk
Bt8jTIcfsLfyEIFiVCQlu7DhSmbcX2FxaSYcwWOGj3RiZ25x4edqHcSkx949mevxF4sEHBB2lCo2
6Ao/3k2ude+mTFOFL8lwNFvniAlaeh/Q5tzpgOoOESZf6xrTJQQ27og/ftVRd2s0Hg1jSQ4A5jAe
iNA+mEQw6xKnqJdpFhG3V4IEQt+zGHKgNRIbxpuur9oJxl8ZTN/y43xzSxjyNwrHmeLet21YpIWP
tacEf4/o2bnqHbnv1Y/yqOgHhJ6LwiE8A5BpjbcCF2/MxMrslIQetMKMwM8VHbeW7IKm4uVOkFWW
IA9G1Iau9TdcjLy9jwZsyxsYzk1T06oib9l2Jzt8frwoyfP6EddqMCPRiQC1DW9b+hf+jKI5rqOl
T8cPNLYSB4fbB93qdowtUpM6Ai279T3BOt+HvnSJ/p4dgBStX6yR2B2f2B3Edzqbg7sS2YqlQo5d
ogiopZu3bKsmfFEu7nar/D46gFkAI9m0crxrPA3h2WIgP6j+yVmxlvZ8qikD03qtBJAJK2LtRFhg
DAJP2yfzdcIj081FWRQ59JxXUP6VQdlVQ8nV5wi2q0gkcqTStvnGZ3PWnjuseI3a++hIWS3acfSA
zD2umDn+G9sH+f75HmEpKOQgXzz21MTgekAQCEjNbQE4TFOX1sB/Dx9zXYOLAUG2/C2iWaETgo7i
NBGsl8VXNYuGwvq+7iUn4hwDGHok9WRhTM1HNdJoa6J34pZPUL3o7mu+49ecrTOlkCgCDSF7VvuA
x9SJY6DfQbhL1F2PS0LSUSplfrhdfZdyJMD2yFMHEeiPedjw36ANQRYdMudYIrZyAtiQRLZberDI
B0q+o9OgoeqYkkFiTN9neCqZ9opG+V1990wNUlL1PZxpXXVx0citeCznlFAPtaMfC46YiPy/Xcyc
uRU74vFmVNZiT8EsSdeoS0/v9ZFgSguidLNAi8EH/WWFNOOBply+B9bwGsiWkxSto+h+IyXVIXyg
0uDx1iKkA9VqmvoCrrFcOcqwzUltHpwNbprTCUw3XGB9SL1LAsQ9FGtCWP9vDPM5pbQHjetCLjc4
fj8+cavrgHu9bFM9Kt9n7VcP1CuvQ7tek1UhHzRlxa2kj3snbTWBpGUwsVMInBgxSeghjCvV0vBl
Aj5Tabaf8UZVSYUDrPVHaOiMqU8DrYED0pokU6Vn2pbkL1hhinU0TkH7s8Oy65GiD4Sk7q61dtQn
/XONCvpzj5qOZdijAuGZs0Bfw5JzXyPKdkrueueC6ZqotcAdu318zo3z8ImdMfmA/mOCWZbIDl7M
gIAsyDUo2WZ2lZAgBErdllaxEv1cunzAkYIDZ7vzwpSw91fQKleGVFZZvJVajjM5d55X+sG2y8ly
kD4O01pbntdOhJ281ey1dVIB5czhR6DRNWnOqFaSnaCRJHlo6S6DSicMoicaJ8fLAJWFUbTGog1w
Sir8TTFHo8INh+yH7oEbnReuKtMMoD0Rak6jB57ne5RvFmjTywFJ7M3+7maCLY1wPpD28LebaaIL
PhlHxjNPWVbugOYy8ot4IxhfjGFVePxzI0so5gcSWg1PRsK/i3EfQ3ZT8mhMs3jRXIS8d8JN+jV0
0KZAItFXf7jepd3llaZTt0nQW6RuYyaVmUCLLcQsRRa1Pkb3XUGt2W3pszFyFCoMc4PuQUbeUT93
iLspvlzFr/BnkgGLTywweW9/6/0EyI6cV5jkVLEIcs5Nasw7AQ7wxvPiciTbvEhUGBqO62YUshmN
MChSFrstywpy4xSpBvZ4Q7lvJJZrUhkSWc7htCblaO2X55jfJVejw+DeXVAKgf5++BoplIi3Fa9+
vmxezA8zP/lWxl5iNx3qZfy5+U6HY3LSOKwMG3Usd5j9aV5ia8JjsvS5spAUKg5HiRU1KVHJmYT9
3qiSckuTrBxw+8yVILKWg1dX4tpEwxIJt/S1Pyi0LAaEs6235GQGtU9xX5eMThl5vY68KseAoRMb
mawSBm1GeCptA0XZ2SX9CtP2HoBF/FYdK5zijJmmIYJuV36/hJnLBFRhzewHVwtwE57H1obRgJwK
4nIpmiVIxSWTyu2qM6Ze2b9A7+9zrB0CCMN4q8wimL8FYt8X3R4EVdZVAYS/bWajQyN5lF1bAh+J
hCMotwojL5PlpHPYtiQ1U/olUjMLoq3Bs6ikM3baC4wm9o4arobCtgfl4g91+JgyPhnD9BUhPsDC
VdMuRKTCGmwyamuDd0Fwu6E74HgG1U1GHWYEKlCL38Ozn/MdDJ6Ak9+/ldLSR4bsdps4fEILMOlP
8wq6fRloxzkX7t4Xgu3QnHxF+c73iYt23c4stfZn5+YA4ze4vUDAONHMaL0/WZ5mvK/USG0pVosx
OGPaMRqRH+3wfTNWNgpLyHXKX6eS9K7yHGorFhpH9dOejP+w3uZ7FHDWPSO1LJMSL+SSxKbZAKYl
ZZ/NpZITdiuZ3wmR3XddbjSwFZKovfNE8aygaVc2JMm4S0ohWhrdRYBe8RtNxOkuhb5+5pmh0Bmq
NJYrr+BGIoj92CvDwjwkPyoEh4x/LX4rSZ8x7PrDoX9H2LllwvMWtpxC2YhwEfbHzKvN+eZ6GwCD
4aOXiozyQRPtFEA+Keku5SSoeGxfFA62TWKoyywmxIg+A+hVYsp598lFSBw9gEb0LxtSwSPJBJTM
4Ah1CTemCC7y1tA1GuGAYsFniSRAIjSIvXYSSoF5WRl7snLPZ0F4O3n5NTC+Pw6ASUwSRwqWH5+1
T7fKVtmOwdctiMuKAIxUhjwHGic06FfDozG2l7Du5Hel7WKvBlCPu51vGbLdLM7YyyRf79Bs4ohN
pWG5SbdEjOkUMxSrevVbTOwdWo/3amIoVdgTH2rrEZhmN61MD6gSVxJhqAD+WzXPLYSDN1nliEsq
V7bh3ELNn18VI1MenJQBXumH/DygE09FTZweIdxkYhav4M8SVKJHwsN9HSBFLqO9XYR3lpaIkoYN
z7H+hIdBTD/1ranfSE6tEuPmPmjih1FeKXmuUfA4iLyUgVIfGDgiRDcUWAxHt++UB0mknf9/mwAn
mG2Aq/sEQn310KVGbXhMtX6p5pUdfcF7OE9f5rS91/uNynxdyQ4aAyQIISxc0ZGwnUsQKD47EXUm
rQfhRVD8ap8G3ZtPyxidG6Uf8iyL76YCifyzbYNB9GGuyNAVuUAcFZmON+WQSv0mljgodEP/RiwU
cqYEVxL9G6tUCpSajqusrc/kXylwhRcU+dYTIvS56jyM56aS4qF046vobpWvh1kq7RfAsuLituhl
OjruLjOd6r0yQ6ATgx+jj9eLWBnlwC/+LqQIFX41bm4+ke0Xs3Hd47KWq1X66UtJL8xk0MYbBMpK
HhOGnyMndW99/vy7mzwwWlO5BzUg7PzzTMNG5MOCl1J7nlpzqX7ZiZW/yUJeD97AT+r06X4202iZ
T9MeWhJVbMZd5iil2f/2H0uTvzSKOWaV750qKmzo5xWaC84SNg17CJ6TYmuO0d/R4sKgvTKxQIEp
xEZFfccUbAP6ZAtATaT2R95R0k6qvDDU3OuDMpjYzEwb30Ttxr8Tz0m1vdL5pM7SFxBv/upSBMtB
k8hJuudHuAqN/KDsJn1Ii6/QzQ2/vtMcaG48FkHeSOTQXQ5ywbhhMR+cHZ9+dB09HQpZLilrQr3t
ZVaB0OAKxBqd00syT/cNxCuXkzqOvmfkpBzTB30UtM7j/IAIob5cm6OqObkH4ejLkVNfggBKzmpf
TnmzkEQ7IBWITJ7rAUw2jMYAkgV8LcQScEFsXvwZLS7f7KeNCTvb3hoS43vNJe9qXzFnAzjydjNl
+wa18fbZRcYyBsnXVienMVG4vzwDeZ/zaYyPQNjg3INaWNLfN/eain8jM3efu1ZPs64g1a77LPQr
NXS2AzfzhQ+9z8xvb6gH+trCX8Sdqt2IoGi9+TyX3wOUmKk3FPl8LyLnpLuPMvuyZ6t3ugzpbYJ3
tZHgY4eKlLuDgb9dq/Id7yHKn3+1JLXe+5bX1G3FaVdky47+j77HT3TNOwZm1nb0M8VjZFA6NCYK
wpQ/Kwjyjrvy7jiLchtgRh7Sw7WFc+kwJO5WjDKrxNRLNugPP0ygiieIrjbtGSdzc/NFs82j+jqN
t/VG7urS3j1Gf3cr5kqBq0W0ExvLh65fRT6pkvFkKgRZKb4h0K3TE7qQMjRLBjsfc9KMRp459qdZ
pF4hY03yJzbhenGu4R4SDXWZUlWtbMDJqq00GPm0KBUzIhbRPQ1H+cl2xQGuuNnEaRNlw+BQRSji
tawxi4UIKwjh22KJBrjVpGXoYaFTIcZvumJdZtcN74K3FUrPUoimGTG5IJipxqvCzsE7k+q36Db5
dLSEdHCk/QJQDEkl0D5bQuSrhoz9/GVbnwiPEv2jKVg9jbMVxpkpf1smqk7G7BX+jNVqH/N9gc2L
hg8W3sMVFMVI/K9E0apsUeyc/XPQBfOq3XnrF9VECn/vRQDHJ0ppO4p6x4vPkzPGO2uvkAUEXeow
0UPq/hLPEEHbhGYKBf2l+Bo/TlgiWDo18U/bGUfmybb8kC3+f2qH/q/uplCjp2DpBcWt+2Mh028b
YVCvcHKZHRbhRD4xNCSD4UG4bQ4PuZSWIzxV0VJtjeoMJEiEIo2NZQ8NuJ7f4C6Vf8Ps/qohZ0Cg
zPaaCFehCMEXePftYey2liWOLbCv8CFjAN6vy6Bj+LD92HJlOFNP0F6LhoC8fIGsQG8JXZ/CHKw4
QJTlnMJByUN0tRUxQDehIBpTg0axFJDLNbSdmvrwIQZRHE6VDaRotdq5sMIT/Kt5lN3OJus2If7Z
O6xvfuXvor1MSCZUroW/m0/iH4d+cH/l68XeYr+3QprtQzMRHzyRltqM73i/pvdxRwhWQro2I4V/
1dsscR/sSMgtQ60gUgHzSLws7He0KlgXPPG6wrqy6UxtDROJRAjGjHSdy3ohmtPW0EycZUyAtmtf
2/GYFP3QpTs7fgRyElfcMm4Go5K2MvRzKFYA+o/U2MBtSU7wdImDpQ0e3Vh/2X6QQRQlyj3p0nxv
hGeItGS49hfqiM/HcirutRnZJ8P8qx6m2b64Jk1YA1DfMs9TDseqmNewy8imQTemUIVK8O5EUmtH
sHcxYsYPCjXCK7iH0XTopjDCQMQJ8RzKIh2K/hOLH7Bq70d2YdUpk7y9Ow2G9EZd/A/Hh+Tap5WA
0CdVmWsBPpt2qw8JGZIvF+hWzyqUWDHYFLA6soQOkhSNbpypav0jRlUD/3q6hBaMsswhDQ2DVMme
F3jPf5rY6wvh87XJO/lICk4Bxwvg5/P9RcMO4FcIvMWgCUbCki1p9Y9oLAhPW24tUd3bv/vmvtpp
98tmtccQZXXTwpwkZJ+/BamB8X0N+voJrab55AQoDivj/0xaikUJYYLPS2JNsDXtYHXd+1pXONTo
y7vJgcrTCszGZ2JgWqRtdNIqK16pB4PcfWd+Bi+WzhHgZPPvvuZ2aTx0tJs42j3UAxnO3m83r1Qu
O8rUkT37ES7Wu2X8KU+UVepj2qYxKzB1KW7aVDclGyMonfLXcDMBUH6LbhlkLBIERuKjS8qP81ZP
uD/d59YFJOKsAzbc8OLLYbkO2OJQZDYAQDF/okmQgXeEqPw9uAYEbnEyce2emRy1iZcD4v7GgtRp
7OPlFR24no1LPOH/2XuqdQKfTcZ/lRH3GrmFUWFFsFXDQJKAdxEZafrzasU2MtVJcvobXy9g7J0a
6CUAWzXjON0hCiYqIwX1zsmuPJXkpbRShn7v5Mu8UxrQcFc5hpesMIz1Vp9oAZCFSAqPUgudfklc
xfHTwY/cnLA6Na2W2iu108v2eNZUMon0znxwe1VbhDrX7oWCIF3RLqe/BcHN8oL6hlnnu4aL2h4z
YUhbJ06wy5qjV63WjEcIn3p8FlL13pHhLtaNDs8ci2a2+lgKzK6QVBCqWzQZKGYeQMFMVwDsZKsB
eTlzHeR/pxM83UVYeb92nCrLTXr9DfJ6I8wH8Bp0o0vSzY/FgfkywqS41mvcTHggGlcLhpSrI/x7
lubugnK7bdKBvTJWOiL9E/yzmyszGYYNvrqsl94QqyJzWt1EwNCOq80vSDsG5oKFigJR+io8wsnS
GBz3of6Eq7T9NnC3l8ny8hhYXbqYG9iZKyQfgIb6NprH2STrPjfmaFDoPNYRpY81cy7kKTsuFAdf
3v5w/9hatQzZboLGRL3RuEo4ug2tswLLkPSGs9+j5p9YOFVi6BXdzpOvjYjYYeEZXTjLZkeRfmKq
knq0tc63WkL2z/dVltD25m8dr9ncSBUJTM6lNhQDAlXe2qmZWkzfwgArcbtLei+3pMG4cCn0+Ekn
PTVKQfSHJUv7FsDaZ84IjiHc9flze410ziBPEz4iJ6WGla2mOb+qd7nN41d2XeSU2beZJITM0cF0
MU3ehLQYFtsDxbNIZdb0brsgkwiviKim3JfN7uQRO7M9s5yor0YkWTN+b5LRxOGt2o/qFos8qe/6
cXXnxKoX5eeIDJBEV5s1+7EDU5NBIbSONuapfVp3Sc57H+0M8wfCZChuVnhOUqT97M1tcIK8I36O
NttuSEq7qxcJVggfCYTDB9fVMLBE2vf4UWSjVj0pmAyFozkxd2cSWWWSIUSWSurYiYibLzJMSHgh
nc6wXh+dM/cAY5m3ZDSllFMTNRzxD1gI1yfV0iTgrDSNN3n136VuDnuuAS/8es7bYJxExRQaQSSY
dtzZMtwSIELzDI8kW/+dzLBwWxZfnPxl01Nf1q0G83Tv4PMSMJ+vbyysKoF519giqIYsuRMYVRi9
MpAKbsGmPTXXiGInuaiFI6l/nqBB/SCuqV52h3euRWoeaDCn7YuPdEahH6JIe1YS9qM2fI8BYMUn
2+kildHhtHwpVi5sl/yF4gOrwQ0npvKze+bkqRyUgtCKfbIee9UWFNcrlHix9kcW0tSiJ4Rhioa4
dptQlAlB4+ZWYOP3cNM8mn+ISmwiPLt3Ds/DMdc5DCzAfMO9gRRL8VsBUjArBBJzO9YBaLy72LgM
JuhtZIYNl6CGvygyvMj69cQtaCRfdHPl0TttMFDsFxCg4Fx6M9GbgDv1Fuf7+x8CBBEW1AP5aMgm
W81+h/8KbgKy2VZU0ykFt+DvM33HTeRp8ScV9rQCaKJozKvnY0Kd0YRyNeP12nkyiRDleYuFgP1E
SyoOueo+EABQTxQK7wx1pD/WvTIMRXNeAFDO5DjtzjeMYU8k7BOOFNDLhUwW8fNqrQqsBgRO5hRZ
YsIO2aSi+oen1QKWWbS1pjPcCPxDby8w4YjKlrc6jo6C4ASNz/OnQkbBv/AzdFID1q+X+arvLNqD
QLOHTCbEdz7fFaGtKCzr4o6e+YpKN/tBFhNHhH8Qfu5llEBTZCAcR7MzbgR+/DPcFWQJ2Tni2KFS
9a+LGOL8XcXsFshZjmfWTyHqsmTA7IOsyd2n885POfDIUz9cAlUmW3ZF6PKn/0nXG7XcaITmQaeW
eKG4gcAIZVB/W6cFA3p0KWeM6uJRf/6I04846avU65J3dU33W4XSeKau+AFqFSNTAe1nZFWsqgpL
YpJnGQKNRaQ4Rt6Ui0HSVsLE6Quhl7V04qet75WsQ1EK23fIYJHOUp7nkVpsnYqqnjW/mAP1uXhP
AFchjUtCY0bp4T3Q5H70D9jYoDz6wW/U6IxhLiXKhLoPdKyYlRQS8Z7u+2rdsF58dnErSd/IgSsD
K8rN7SNS1JCE5IBMH/gQabSWts0arijNRhYHFNWkGEygHG5En1mIqZsu7zijcPDJ8trvVWj7U2ye
JQZKz/AB+IlzIPlCiyODWCZnQgIoY3S65wQ2MF+Czw/IWvrw07l6toXakPjPhWPuJ3lcwe5naVHW
VuNV52HLFw7xJYYTl0MDeDENsHPl02xTFARgIrhFtwEnLjHz9dd3+IT30YKlAxCmzM5XC3W8phHF
cn2yoqfeu5xqripM2dwiEJPQ49+xWYVy5eQv8f0QP/iKG8tLttfTx0Ok9TBI68hflhytFDdsBW1P
ey69sr6b9rKuhezlCrjwFHtsfon0qQPvlljm3fskYiyvXVoTznSWr9PZiwt9wTcj5XqYzQAxnefP
sWdN4Dz7hkBhO/eH1QmiaLbBwF+SYs5STmHttbgRUKmWIkK4XbXJplbinmXQTr68YF1qheR/ZfJJ
idsYquTk0RX3LjqrFmC/QpWJuNKvXBFm3U/u6EGS5wSZM3NSWvH/Cw2b+Acna/M3vPsRH4GTcRZH
Hdd8wLgd2YapqRdJY+CQlTBIp1WIvx8vc/dib9w+E4+T3cV87MPTg3e6b3du+pBx2emIkhlbg/6M
MDaKvs1b1nGD/HQNhYJg/YZWv96JRQEb0iQZ0ZPje4SsRF41WiXBT+PQ1F6yabC3NEk/M4emKgEe
Fr6pj54R636cMNdmd2xQNflzsJ07zqa+G72TdkXvUwtrkMxmFC7LURSpRFU365WhxabVgjtp4N2a
5SWkoKSRPf38VxSTKSzC8AVLjQPgkmp6J+D0hcunOHEOlHaz+42CH/g3fk+DMbbMIRKKtbnpTGlP
R22wnabGirJKS12LEvjraVNCpZzfMgq2Aus3QvmHbj9ZepK0rR7xPEjsCNlFlgdzB04Hq6BEQk3l
nYUvH85wITDGxHzjBu3p5ua4939fVCkKC4BIkciKmew0D8J0e68qsF1qqDO2zJtSTky1WtdQ3sUJ
Xflopgt3SEo/CRcBnueoQAJ0+dotzHAgNXB7Zd1Ii6phqyNja1w/S7g8Bu/YQBLgeREdrGQFUw90
f8P6LVYPS+n6J438+fHo0/0y/INVYtXdRHx8KMH0lnkNYkvFtfEh24vsCgVRDaWzO/5nAi+rV7Te
xgBM3UxPxBguv7qg9dyHfDXH/ehXNpGTMi2gITqmzRaGiWuadB5pnanTcpkEgrMpBXuZFUOrmzK0
K/yYhv4fJxoHw3RbIx/GoOKybv704NZredeL2ugGvVO8A3RiTHgjQG8Vl8ARjVVa01Gd8COU3YP/
TUIJfpLmh0hOpCVRqTKZUjQ0FMVed3y5C47LxSJVGE5XG3/OnUYrSoBMzL17DXXprc2a7/nbmkft
uU1wAK3DD6I5g+ySMpaeRJ8o5jpyQj1dHmPvTkWObnz+PjkcmnZ7UMzTUSnrLlueA2KCdD9V0DZn
t9ba6s9f2Sut2p0WyVk2UH8rBcGcOu8oDtKpqmh9XYOyY6mzXbLja6EWznrg/08QVSP4bnwULc8s
Tp175Xic2trapHu3vsnMxCi/TmNIhX3MmIo4g+4xOdE8dHtsR1fp2MSFmHwYWnjT3WLQax2LdbXW
FSgu6yCfViaZ25IjHb60I1YOBBQP45KE11WfVCUndRegU0pKwlR+pDogJa+rM465VAsqki/ogLRu
Yhw3TJw4LAFautqgO6zzki3En83wfZqReAyFE2yR3sJLc+QPkC7ab2+FU8Cz//PWU8glFMDoY/zM
geIM2NcFRo8JHpnmtF4HV7Yo0aKH/xcKFmMruhedDd7ezrH9q0XEbdtWN18V16YdkvRoXBDVQOXZ
kKgQNKRX+DJPqneBu2P6jtrn2Q/xQX9ebDyFryNw0fi0UMXfcCivLIiC1be9YBVDBFkkofO21ey2
YEPHlnbgxeiZ0qv/Nt8OOyH40fCWrnXOJSxdoC3nFEZgf3dtfu8geUE2LSyOCbMlIz+mAGg2BjDj
ReGpU0/ChVBN//CH8MnpaQO/sGDG/qniq/0O6e+IBuFKuyT9bd7qu4tGHkVqy30bXKbKpXMWchsi
prSNhGlaWHZ8Pwe0G4FG8WLbcrnh5rfoDYlWxTcJyd1BYZrTyjhiPtcfJ+8Ek4Vp+DTJCOgqtETL
y0cV9X7cFlPIOcy8lSwRYwrjGRU9cVUfUKR4Sx8UID9EAKqBKTVSoANZTj+fpqerRwL8u/5cZR6J
cj9NnB6mtunAff/eUIZxrKlytRXDHgfkU20MncP4l2gx1KfFCtNKFTrqpAm1laanXMsG+WJxWAuB
J10R/5fgv5pPly2GaQoRqCclA7IZfTyAQK6GNCD1QLYvRy39Wj9LpvL3VeNrvplqXUEqCElCt35t
4A5x1PM2/wuxAmb7VNAFdTwBeyA8YIdm3jA5zV4oqLgib3bGfb50yFUtA4reg94jgjpHNkjzPbS7
nWZfsrEDCPDdRIJ1i2CwLEKuqMJLISdgk3sxZjnSz+E1qSUc/Vr03aWErp0dHosVk8IJv79Zozaw
640xrjq72kF3FZKFJZ8w/Ukcnyo0KvAu7ooHis4Qq7JgSsAHufMLI2X8ygC+zZJ/8wPbAiVANKSn
9Yp1GNre0fxUzpa/g0niHsWgajOUSpalWZ8SYW0HZBI75Piz2e0Qv7T01jnBkkr/daXsUEoZQux9
uYwo90s3lwrxuuHBFiegFAl2SP1jn5F/RGwjm7W2PUeZpSyJaUDYDRwBCzvp+djgYsM0jxXKKMDd
/P4u6AeWhCIFTYJykjfouz6x5Wn3Uiako21gC6b3QD1whr2eXJYcnC6NuzmICTgutm8B/xlQHe1e
3KK1oCbpeZdAoKtttI2RbOn/6Ot0DInQ3Nlejp6AHEFEPoZWmThd1u9AjX0Kbqi+dOHAgI7R4qM7
HyrL3gQFNIA9xio1/YOk/EbOoNdtTjz8QMPbta4yhddGMJTtTiq3+7ljcgqDNaXlHit2Q/GcgyRE
pFoJOJd6Ny3uHT9rCwrxV6DcfsABuoHp9JlTGSVfbM9Ky0/2JsZjOef5KfuMz4aVCYXv8AWHRDiU
b3MHb2Xqkfv+dZLedyktGGGrQBIi9V71Zp21pO1XQKBFfyfVjv2/bsOTCAOtB2I8kcIx0i9ZYwLb
bWsmV8UapwmlBqTDnB8SRctGi83S1pZkiVTWfROTb1BVXkAqYopxMQQssbK9012XgSefC8V+rXLl
fOugMHFQAFMDV4rSt0LvGn1XZS+73qw5cV7ckDTCfNEBqAHn6D2u0BPIywIoBAthfG7auQ/VxCIW
v/2HPiBZ0ELkvCdH/mujE/msZumKoQcP/rwPuD4UrdERNIYibpf21RSh4gWJaY4Po/hyxard/E3P
0Pl38CI9jy8fNkR4tVklLeGOyvnPFSqx7d0nl0AxKDEvQ4cVkI5iNSsGNn8EiP+ZK9OdbQoW9KPM
bGDLfuCJd28AeIelRjFovZF0FG+PvAamDQylaTjZQAm7pmQcYUPUtOiosZ8qDXV0THOyveGoDurC
p36i7p5BLE1XekjbzKgxCx3BD5IYjSszL3Xouqhgwq7uFZUtFM6CpZgVLzUoNfcDuTaK9plA1VRH
IbDsBK5zClg2M8J+GLzNhfkveXucn5FUE5Ii0bKOTObejs6pxVNso3oiH51DkjlJowQU7Bbp/SGK
Fy/KmRflYYdwdLNi6eMmOx58qWUn8Y6k4amQPHUNe+0d65wBeavVc2ar9whZiUvJvlsLN0AauphS
U2ymIzXNmUcEKjYGoRxGqFpnlkEFwLeX8bo7HMHZ1gSpRgzDmdv8TV4dXVNfzLD7fEykqUdCgxkP
FktP2TljomH0Z8sou9sesCGSScCA1VaEhDllSsJW0UCyRBA1acX26TwfYCnE4CJzljkR73G6wWjH
mDTaGhH88FAXYs1jzgbKeQs8nYRh1QRVs6MWmr/FojJnz36NfLfJSQSQvIb7HsMmxIxwBJIMrLDN
HaJK7m9ktzQgm8s1P5Zb6DGHhwwibQOFyvHkYXfMIsCsjyr4gDzko6cJkif5pFnyYmToi8Zvhixg
glorYnEJh1eroPPwBwCOJyf4IOfWrt5mI/pWbvhUh0W7uChwUV7UNTvfIQTmVNUj5u9L4t23q457
65reBwZdKM03Agk78OsHxoHq89GiToJhmBwq0/NMrkeTa0O0cyBaH1u7obQDQ8//kURzZjA78rNe
ps102uLfDR/iGsm1DB0y5FEyk91C6uIY2xiLgcGyQs7b6EBhBK9oRHnZyN05pZPh15L5tbNY+wCX
3J6YcDbcjLwSswQ2FTyYjmWDeGdpL5AXpanCacxKK0UPp78E/QVHPQpd+w7i5psvNMzW6FjeUig8
FxHRSNm44kt9MUX5xz9cj+MOkaxmqIiuerdA2cAuHCUi8rvipPPPLja7Zv92WCNQnxidBsF1VND0
uPmPPzmFBBhsFmr+bWMOZ8zzQ+bmXaKyEmefNQF86a40pE7C9zIkBSrFXDbp0orU/n1wg6IHzMVY
Fk6V8sTD5kBByQX0fugSTNoyuR4iGUlMC0SEiwuFzNAbO0bU3dQ3c4ZqA63NPeWbFlq0F3aKi6OB
VMjzm2rBhxRJTl0pVKsM5go1vTLsJ3oXn1YXtVSRK6q9OpfAAgolrw7ejUtluDoxOUtLZ2sNryHo
r0zrGe6P+B5jAD33hkGJSLgvcoQSkStZPkif35yWdAuQgq/Pb3+AUoezyEptfq4q1a5uBAqUs59L
AvksBzYO8rOR2b28uy4WbTqCXhQzpJKz/QbGt21+104aCl/+aPcifWB6k8kx/OP9pTAvPVRiJdNA
xamJqH9Ktk+8tQuTPQzJ21FuErYNJVWdOIL3Y7fjgrQ7oLjuL/LsALUoAGMK+j2wDhG/SpFT0VNL
7n/S661p0vZ7hqzxTDHdyNNH2ux1kj3vi4L3jrkWZiHlriyT7zojjhoXDuAstuQRxe3hcFNIW36Z
Q7uUTxMstgZN1tKOytvfBwHBeb6y6YIoWCDRUOKM3MTpIPzyukYHDr2A98vnJWYfIC+DTa+BR3t0
zxYYRnr8LAlWihtWTMV8njWPYRyy0pp99vQw02t5c4GW6Foht0ReQFHHZYp3a/DpIQa707u57Jm5
A7y7J7ZQcDTTVDXVA87RGeys2QTLXNcMn/6TVokTwXylSjJ5UHg87s8WXAr3FB18MkK2s3Pzgp10
xZT19iMWIoxGn0QdPORjllCDNDLAfNDpiUEbqI5mHDf+zum1ade6bXq8eVIMJjMIm7sgGcOzGdNp
W1ffed6UeDCVFkeU/eIERO7yncgG9ZcozpnniMu+Q07SosiIxHy/+gqm8ed6QaGsNbVOY2VKwVAG
vSUs4wJT/UEM5HLUCWeICX/6JBASObJfUrpThFTTlMX5la3AnB+KCrFrZMEoc07MP/fydh97rTWn
W8VQx9QyFkqJRriPGNZ4gAY9Eb6Y0Kyh1WhyJXfoCZzW6spaI3Oviu6wnOaK458NpYQ0HqHLrNtS
2Qjjjgu7MjlzVSA2eZgbizX+FZrFcZ1IahzVWEcnrcT7pDFGMLuLj/DAIeXpPo/5cpybJFBpMoc+
PTJIQFI3ehU4w3aNHt3leFQph+F3SIkf+asbDtitzg4WNhOCEAe2Tr09e9qc2UIBQlLshDniyeiN
pbCZO3XpPbVJPgA5d/xGc9G8i1Bt7S4+s+TdStFFC53s4ootXKTI/QrabDyUgVk5Ct77goVk2Rhh
5U8TSJkBW+us6TAmBv/xVJIYLzBcJrIsiKzFYqh9tkYiuY05D0VryvkEZK8uZ3ghYfZmqhKSW/xP
HoGHyDU2R+VyH324Vofcme7I+u5lTorqJP+ORkuadR5nnWQBEjt0W9FHh/365+7NG8gbje+iC4BT
d6K4WRMQWOf0ThurZUexEC4h+MPlwSVKiSPSYfjh38Rwq81EgiwWCiWPD1IZkPoZaFNmekM3LxwS
B1x9S/OclXev6B8sLvdgHSbLZrfHxIDZS087OVRIO4+BbLhbJsHNulUCpU2iy91xdHNTNmDt19WK
2tYQuKs7QFnNZ2DhfQAkX1qBbve7U0bDkhQigtZgbr/RWpFREaGbRLN2Bv5WvylwKwDnKo8fgsyG
Pajzb4xNV+8mmU6H9rtgGt00G/9Nr6tKto+QQztOXoHTH0Ttx+rru/HIksYMQP7K3XYwm7uW2Ige
sRYnB7N+Npf1XxFUlAe3/6I0oI07gGqZ4Rd8w2U16fXv6dlsWIa+6ZpbIKIC2SdO1LewVWcmx2Ot
sc4zvGHcfzhu7sv9QBzRPTO5J4gH1qfCnQ5ETarSyVPObgUF6rElk0IxtkgNqiO0bAGWyG1uw+AJ
nMhVdpJtCzuS4qp4OAwgzqsD+xG6t+ktQLzJGDCIHFENxsaSkOyDUgiKZQgLkWMi07Q5tRHKdoTC
O85h+bs2EmVZLfTqX33DzVVAdvdkQ9B3fjY3ylRcM2Y9FeNPZ6DK2lqnpFxH6Ob0XEkmacLknRZG
c2t5ES1YVsumGu1uZ4nfV+3yDOt3za2geVXRSh3LSsU500yS3NRZaxYOYtn4ku5ByXq9MF2kmfUw
QWu0G+pRrkYYADcq8oleOJHHfSyTMt95pWErj4GlGDoY7tZPTuBIsbIwoXxCuqB4NQ+SOfQMfKmj
cPgQUHrrmmZ6jg9sqFY8uqx0YYWBT66lwALys3WYhmhthx2M5+32xKZQSoibS7tMUUV51pkYP6xb
LRIypjRGRSTikLXsJkDimYCeDoFgYDSy+WfqKg7SL1l0KS5Uf8bOMayrE6D1eDXAuWl4nZSMUntg
EBhNpfbu/UWDrQ6oedvpLDo/DSEA6/LtRn+wHmi4xgV6LecP1xhnQNLLeyOzm6alHXUFauD4XyXX
oCphD1p5UrNb1sv+CZ+7TyE1uPb1a0zn5EiVkbvHQvPrMyYVu8lLu6VfWPwyhLJqtEq7UwrEoC4S
KvW/NU5rtjIv3rKOSzPM9XQ1zzK4EsGWnQwomcw7rlv8X5HeO0YY5Rhrm16g0ZcLpULQYLTskG3I
mU9Cll7KppY0zY6La1v8GIm+WoT/1S71JXnWrIEXzC/R64P7SHXygrng63BzQSmyeWz8jkbPC7e/
+MZQN1EoCqIeApQW6oT3uKtALLIgOq7A73Mq1bnCf9DpXTniE0pReEhbTP7IuuOxnWeBnySU9+lU
I/TUP9AWtMDG0JCq+98uyxPj8JWRV/wO7tDQxlXwNaHHVUiN39Jg8Ai4KHRtMXVEogsxpyKWxf8m
kBGN1IYpiwCKZPbEMxJY1n/mwHc+1d41AqkVZ3V1F+4AC0BOH9uhacCUe7xdPJJWtS1YKwHwlIal
n+RCG0SxZxdXeX7sz4scK+1OmStFGSBMnU8ghH0CabHoHxyosQr8JkprefgDAyRoKkv0CnUkPYFO
TKtuOs3fjTWMUnz1EceoUVsPkOPh1FCNxiqitZagAVzRod6iMinyrnmUg3JQHCp85vIioL++4FL+
tpmzf3OEZ4wa2ifPQN8jR1N0INpImCLQIlv4FOVy665PUKY84i0nw+Vb7hb0FRSFVjIRGsilB0dx
9E33UydF3k0xRl5RdMtWHljhLrHhzh5UTkSfKpZGAn3NSUzz8cfRFOLd2g4vWeXxlGkch/7ubHl6
i72Bts46ohhL3Azd7O6klfmZxxTCRSf7ldFfc1xFueqtApjtUGc0YZh51Yeuj/y3XdCmwarvxqgF
7RXIleJqLUeBfc6TYz8q4ygFiYfWYdQAHjKqwhN2MU/PjODRpa/kNfbDfnozczCHvGOGi9FqYgUi
C78tqjz2aZHJDafJTlE8nbY3A/ajXoJmss+HtGebua+g1JXHvG+OvFhmIJoadSgqtTmN2CWRuD4E
mrko+BQIbcPB+b3KFWTjS16jMLo+nfOgH+j1463g9PUxu7vqaDRD+GUhmKG8dGUOoGpgaf5azq9Y
wsLzEfzSRNQfTB3KvQ9vlIheCZcErGZgitlMO8fxg1G3FQ4jmBFQw44e1l8OjHXLAqWv8o5F0dIr
YKKbsbwJLz8trPHlGFwj/ChMkvwfDaUd0DegJf+sqEMpG2ne8LrYzxKpe1HaIrzJoOZcX24ONnvq
lyHEjZWk2jZW3M7rrBC26ImGf3d/p/1OusEDrb5VWqcxUMQB0lmqrEtX5LnhoRW/WHR9+ZyokguT
Ohokq+X6CYsxeCO0Uwnwsmy7/EvZp1yJaH7PWP5LTuXOPorgTvex0gsdBHbX8E9/+Lm9SDEo4ynR
0RYtSR4iIERc48utDxU3k/xEgkEv5MDvtL65cb34bNsfMTynM6+MUTJM5nxMjNJwiacWQiFaL54l
V/yTD/Xunh1Nq/78d5/TwoYC0UU8ZftWYrJGQxBj6NhTeO8CGg0IV1qvcG4bje619z0lLcOmpHj4
0d3FQOAysbCwiIdjzSu+MoDjhAm3PFMMuaHdqulG7ZBC0x/shrH1P4hfqt/UrarF/7MYlV8wu75n
Dc6e+SGpNjmitHwQUZhaFiRVkpSpC+9g+qR2XBlbGBz+XvyWfpkOHKvYSdU1DDO9O4uyXhA9AljS
U+FKXKKSlCWwkV6wxvI5Ldx49vxahkM1OVg+cTWUTSSnV6BCsNCrQfi17qgxRxiPX5VNPlZ+FwXd
vv32C4fuaSC4Mzfnkn+rW17CmdY1Vj1B2Ta8E4pm3FuIkmdXN5Ie9Fv4IYlYtr0sn/2adYaSzMwJ
OiSreS/z0hbqrkfrZ9jILu+CoBMV3np4txUAJEIu4lAwcWNwEalfraGGc0hpMuIsV4oEKJBN6Z4L
7t6ox47hMqH0+EW3cloM+ruaCnXGuHq3YGv3aEepGRXVeNYsyC71Pn84yNcBLGv2TeZjO70s7LWD
921CFwIStNRNA3tBRSvKhG8UsDRNgbxoIgxz7sJH5F97EaXo1TdCbpCw4yw/0TYbCTScpKc17wli
MYuAemGO/jVZmpQiZVcqTm1TuU8OCQIzk8Myt14DvV4oKaLYVnGr/4tXIODQ/DOHH6QAbVSEN5Ru
DraePNttQZw37gEFk7y32YpdpNd9cxxeKaURszOLPv6OYNrKlfGorG0gep+0WDkuosuaB6pLfvQ1
mgbOpbVsUEsuwZyk1TLYBR3WeINX7CHBdHytP6KBeEbxZrEKwnmQEQhpVDhW/esgmAH6wSJ9prhq
5E2s1HLnSgZlMqjRJD43Logh1nRoHFLVCToZx8H1LADw7Zr+OtDgS6F8Fryeocir+zd5Fu6lynqf
mQ4DvfHiDR9KuqjqHWAB97gi5OhutzINtOVXFjJuX+1PVxoYJDqDxPuk9grkpZLDPGhBAh74/aml
RvLFYwZEoSSbP9xwH5BE+eJt8Qmb7FQTQ8gojdLsjp51PMbgrg6iAHUCsESBdY/AIYpmTWIBflnd
SqYUPWt56OYXtyOERTAcClLF9USZEJG8tJDjp/N6fF+1uDC5vtN7RP+kg9BBlsOq9g4UvzRFRVJM
WLMSGbYbFPsFFhjOr2hfYkgt7eNGiXkulGsyZSrtlL8p+zLfE5AjAsSz2IPrNqelrwPmX+g+0GhZ
dn9iLVThMLnOEdAmIv+ncdxJG3bLXsKpvWBX0Nm0QYGFqVsLfVso9NnEwVBqFJbUs3NhIiFeW4Xh
iJb2EIi7xHSxgG0/qCZpeJveI1Kv1J2k1bz7s6jAfOfn2WgA1KY3LptvrMjllbVqefEXhJNfXWVC
n1wli7MZTLzgexvMvVZE7IRL4SUyLH1UZZuORf3/W8Y8KscaQvqL4JuXk7R1gusruBtNfgU64VcA
UsjA4IWEpR7DvOIfznsI6K2J+Yej18dwivVDuxFBbcu2NGL4xZwfl6CqQ8w0QK09sfqs3lGHAO5v
oS74Wk3nUWmkK+Rmxr55fOsrlUECKuMWAN41L7ZacRRIZvQ1oQqwV1qLc9scGJ778WoOSpGgS21A
s7pH9cDWtIlisUusq3oRupgW/Us6QcjBU0ByJCQR6xcO/tMds8Zg2jH7DC7uFGUDGgtr7NjsCxyd
9GIkGwC7L7ChYr2HAvfuwi7KUjqs8FjSfeYfKfLQIJN3202tGhorqkSG/D3A8L0jZOVQBNh5Zi/F
L0xAYvEeXfJT5+7FWp+BBTFAwVSHN8ceYlRV6RCIdwPvL4SFXU/1InJmhigzZ++txH0CyBEEmc06
nPwdpYTVUO/VHKyHWeWWVHpVrAofldLRDWIgeHDtRStA6eVb8ZlZUGKBWSoXPfJla1bh1VGxGhhO
tePcw/DdOZww0gG40DD58gXqjh3olVfmqn3J2AJw1dY9Xn8RMFha2fsy2kyIIf+ZzUUB0qzZfv+O
s3IILlE1Nb2iX7VYkCGV80DR/cwLb8UHYvWES+4/n/iSizN45o/kmXP7GTvQQwmIBHxvVsU5GdUq
0pWRhvoKIlDzI27lmOdZN/2L2x1rNGYPdTiqdkMq8pWypiZ01Z3kYJkX6vxF0IYFa3ZylQA3/O8U
OyeNV5So5oTSNS7pbs9grRuNGjqjz9dctKoqZC4nythOJlxm59Iu9EymzRsjsBkPNM0lqNyk/nY0
oGV4Jv6oucmjl2371+yihHvN4QGjgSGBZ/32nNXPa7qMD2x+ycWYm/55KpnDLn7rg5jb7xYv70zK
oCHjP8fJhcbd/dYRnviOKs4St6egegLciul8V8lD/G1cqH6wQThBk4qUrbMq/qm1/B3mV3XbUuUV
46Ka1SWGn3NtEanxNhDv4ljHpF0gEzhM2d5l8s3Zzt3A9TpMPnMwpEerHuUR84/0+pvKlG/354Bt
V+sUn7M12V/2qLxIdeM1vzsGjJ1P7ptUdWcQUn0n/uKeBKz+RbUe/hO/aQMZ6trpWKDcowWjYP3d
r5DSGKIvZXjMYlhdKaieYNAIfptjUzKI4pOLsonVIqpJxUkls5ucXGHopomfR6fWu/ndVHLEfPvW
T+03WVzc52RNVKfzqkuVfG2zWfDNpxs1Zwwv7ULey9dMS9YJqHOpXLM5qxUfPePW9LOn/5R6fY9h
v/cTeu37WaLWkDen0wm8zm005TF3mxb2ZGzFmlaEODwOR8Dil6szbbhIpnB2WjNL4fGwZd/c9SS/
EA8qTUxDGtMpeEvq6cSkZHMtXACkNqptK50NcXgcgcDukyxkNbcKhX9fndaUdmFUSgvccHN75NSw
ypHccJ4DlNhsH5Nkf7cPkcLLdkgn+xgkcQ/wn0Hpv62o6EAhkhgO9F4/skBXi2BPgGTwTxSs4rbM
hCPkiZVf9MCEiGTk7gI8XP57dGRYDPk0hQrgAr7JIuWkeu/io0GaCzPXCuzmYK1xifttr4txM0kK
jX7XWDms5n6GzU/6h1FztoHBz6K/Qv/yzkFvre3m7AlQS/7+Fu1oxfrNoqS51xvZeaDo8hdtPqR9
Lk/30c/vonC4cYmh3eA56egJHgN8K6T3H4J1eHmV611pb/Nn5H3hvcVhzELciLPc3Fr1Hd+342oI
DsDqKyxcIJ3plHlm6jIhCAnJFjY5BiiUdyai28zOHHDXMsl4DscWlVWu1PJBElYpI+dXPT2Iiwvz
HVdP6ueEkj3EGUzWSJ/laMpU9hZC3Vec0McWi+cSoiP64JnICeEIHFhoEA71w3OgrCjUQG16YwUJ
gXAVpSsz57cDAMTDGikDrCPxMPZ33C6RG2u7kPFjr+ZCgRpxYuMh1Lj6dCfmA+vvTG/jJZXLPplo
Taz46dbS2vLSsutGrRcHdhSRozGjqipR138rYRwcHfiVMhotRer9m3hMB5tDdbNNVXnk/FRKbde1
d+yMXrzItmJT+Ja+C//A2Nnqnz594YbqfSFECXw9X9agaYG8IDLFHUPAWfJa+LBQg9ErMIGGAbsc
w7aVEl8vL2h66KZ0vmnu+3pfv9mfND1xaX8heQVPKwyK+OBpHCOpmBytpg0Ljf9iu+pWlxJgUp3W
6t+E0wugvqkkUuiaiPmosQTirnDM3pEPiuqwKz4ZDkx4meaCjowSC+r33ThVgSBO1xGVGB6cMHdW
CM/tSUcqyOquc9/QsHy/ojDPGdoTC0/oQYzpMNhRBh2OZdLKGkRHWsuck52tsVZhcRN38ulYPEMV
+g98pKVM3vmbexhw64J9cJpwmm2IcKh55ppCyXVMjbFCSSn8NIfvkx30WqSK/zZYHREkk0OfPcqC
zOvnnECp7zW8QKKhRX631LgLDGAaagMuox+sbqLparpZDxL5ale06jtqAZTV1Q7Lx49noWia7PsP
/Az9xQ0wjxVuz6wwVmv2NK3HsdyPx8ufddWeTNyELs0RCRtcHgQQmV059dMMYWo8WL4thBNaFX8b
47Uxut0n6btdoyFJfAEpXLQhPsNIQqMl9IT35HIitCPMkXyLRr4FfHJJFpSp9Wp6k1wmq6HIfV20
HhpUSwEZrnx9Lze6F+OZoZnvga25vg+Ik4OK68DP7K+dVv+N0AqsBUYk+LN9Hbgu7aR/gmDJub01
n3LDtJ8uPIOn+4vqxKECsy0Q/mQTBXt0Q8O2AUOIwihqyh2wUByvKli+CFI3iLLBDzLH9dB8m0A1
go8kVXY1jfpTp0C4o/rfpKcuHaztR6cdLBf866e8di6BFklqDJWGzd08uFlm3JQ+JGmd3W3rJ9rI
Sbthel0paJJj6SP5QQRSYQ0VhA7sDQ9mt97PhIhZKAAQuxj1R4qu+yGzoVMhQCFsEMPA3VVXAVJQ
rzppQOZW4LV9g7Djxb2yqG5ROLYzE7WThBXT0+At2zm7vajBhwexnS0iPQm2NBSR2RhJISyYAiT8
riKMgU+xK89N00Eq+/eaSi7skDqFp7FkCTBizvXsqM1W8iLl7nkmvXRlGRgWphjS+rHnjl1TeeRH
jgvfYDsNaIigsdBJ2RvKzNkOpu4aPjdaLO3t0Bal+mpJ0Hpq1tj3Fwy7h6TqqLfXKI6BEG1iwZC9
91fD5UNW/E9FUu0gYHcC5iCmbzz9g5ec2/zT6uJ3glQpeCl6hOs1gUfGFW341phlIMe8Hx9G6KJQ
aDKmfdDhvAw9Y8tgXY6PlpYNmbQqYAsdAEceoyZLVuX94MGYjiaubzmD7VbscFrW4jwEOswsKrKN
bzhEECK8d0Un77n8JrX1jhXZPT0npKGrd7J2zpam6RY7RxIYRa6hwDubgWwZj4z12S2eSfRXwNMH
cjD+s9JVd+8eNE+wqn8Ae5LHFkrpaMRQesFi5jMkrewVVT7C2BJGb8mpTAi2PZUP8RED7FJC+MeV
fHzfUQJpKUPWn61WLjRVFtLGnX4D2pX55aZA/GVYrqVCtsb5RfUOk16agd3YVFXZxjbjX2oBqHOk
UxXHiWY+QZu6iqfaPjfabc3hPLECamlP0pXyo7yj3SnbUFjHXIFUxG/x4/e8K6dfLgpQlpWGgLgL
Nv+Po9GrHa+rr6jXXkLZBiTBabYgs+uNNh6vbkwxBtNaLgT8+bs/9g6dMgfaq2++OOAowIuBWB0g
3oJu2UkYV3F2XB7H/XIkedy+opnbDKp197zcfYKRKepT9r20MEtVEXOWWM6OREqzlUj3iP+KoCqs
mqeNsEa1dnVImrnhjHIQT8Kh9gy77cIFUeotiSAwYleWUSheeyb+ib/ZoTTjTIID3zti8fYQHehc
7/r4YwQZedc9WMd9l6xCVN4SAo/R73ye+id9/nsIzivs0YUCZIgLDKhMdzF/VH1Kv3RX/uoo1XPX
UmWPHZp7r46fEJrF1nw076cExQMQP481UYUf3FGlTDhjRhCzda35ltHgd+giFNk+qiUumnZT6pIQ
eRA9y5x+qKrjM3x7GnG8o9qICHt7GEseYxhLDLStq/eLDND6h8SEb47bEM02mGszlDsFoilCqhHJ
voNm2+hjQw9eBH7QbaPxZ2uMNw0DiyNcIg5RyAW35gt35a9EMU6XeOKKaK+28uCNqE/E4p8tYD6o
ItgNbpn3XHqHA9BXwJ05d+3MN9UA/cNSEsZs8v7HSmups1qoDmz0GMrlWRZKX9PHElapO8hRZuyN
mKFXBrw/S+LjHYGCQAHCmaCQ+YY586jm7Sm/6fjrr2q5DnzWaQxvFik1ZGrsql4zzGLviQ4WgbAY
Pua2L0PAwM2TcbBA++U4zvwttwz6jCMmkkvqJJ6OjdioTmZK2v8VhDnRiRfGm+3YHUqBTevMjnkU
vqb/KeojQAyWEoSlFYPB+q3+EzeHC3t7ubkiLzucQPWnK2ryH5PFKePiamihaTKygAALbDQlqPfG
gmcKh8ysQLhBWBTaaXtrIBdPW7nsl+f+BKoyORpkSLLdK5CKE0G7C9z53JxBowEdvzftsMVhkZng
gPHG1VrZt3xHbO041bR0gg1H7rnCJG5jFckYyJTAYcAGvH8zjQ/cISTeDm/YZ5WsCNqeZp1Sv1+m
zNEtnlOemsZk0XbIkETxbc28Bl1zGpDqyPUklw3h5BhAxy0DYWJBBvqeh/CnOpPOOH9AceXJlWFa
gakOYAzMs1acajcsfcCW6UbMNBTEM2eLDgxfN4SqAW60hMBJL0zxBxGND6TFrjMqE3uEWGUS+1vX
uVvmD7o+y9NYR8V6Slp2lkrmKRNf5gMk5P1V1L1D2RgDS9tW/E4vaAmLjD+ngyDESOYYoy3oomhw
7tF5DQB++SXAPsQIv3Bd0l8uq6m7rBz/TxpBeanzf1KpnZfs87YP4j4uwfU806CjBSSnel95e4A6
1UKNcJLiVdMILd2a5obRrhObtjSwXkt5v+3i9G38WqZDUfLidHmzJy2nsZVvav0R96JfwhkVcD4e
XVvZ/CxOIZ3G2GrbccDPksfLHEKZJl8bTsm/ERTifxlFDFTTih3BL38zO04EyvKprt96MklwV7ir
OBhTkwRn3eRpVYuH4NGjRbtWv3f0qcdCxFqSD8Oghwox6bJGl7TpIbA1ktWbWhU3DR8bN6pSUEXs
erUhdon9dymertUM/MC3/2s++sk1a1sBEYeqEWef3aHsyJIW1c7S2X+qA1/A0sLOTKztrRBO3z9M
bOBtRAPgbi66qypb2jkP4HugUrmFULiEnB2HAfFBuYpXctqYib2WO3auhYn8QJw+op5EsjJvPPbs
DuSozD1Ux68gJaqz9hovy2enzr5Yn2zi3vxsdRRfsEgQcyUWq4L8T1ILdO9fLIxY+x2SV0027ZlO
HUDeQYvyX7fvt6JIXGQlwsAzADnTdu5flV6/IyCLHcSWzJZYK7sWqtjloxMNKka9TWyxAyrjgypT
dMEbi/K+OVELpKHQsPKFDgJS8FVElc0DIRovBkpsjVrX879eO5ac8McwfsWQeyRKBXLBB28CSsEK
EPNDjUQ/y6GezqnBjmVVGVNPrATMdiIYdl9bp1hk+w6YmVQWAZRl7z/OUe2DryeKzxncDVbWNuch
4Eo+CNgCwMsU4iTBFI+CMCGqnRqmgiylz3G4ULxlCk/ZJS6kEGArMrgtyx1p4Escwsp9uAQ3K5i9
UcdzxPhmZeYHziihFHHPz42IiodrwU9JBhqIWg0/TWLKyfqWqPj08dh3o/wUa/kN2mfs9uDv8zVf
L9ysSg19w/D63dJ3M1ugmOCXwbv4oogeHSaF1XwQIrq9TthJkHZPW2+57IKakkko1EAyo+aBbk31
I4mC0pd3wgCT+Q0Ad8pHATFk6d/zWYzvM5h4F5KOyZc8plYa+N8HQHbLdRrL0sBRfZtq/R2VMZ4w
I8IgwyVMsSxd4m66iUVSL3GjyTskk8XAO1ISTKdfiI8AljiOX5kLJhZPK3SQ9ycIczV5Mqb6Ox3i
G2tkp5FP4LB7oGnG6t/lvmX1aw5GUmBzGX4X4Iguf4/bAJDr47Zzlwm9hmoWw+tp4jagDjkFUWAd
uI53upaGYvcRvxkwjtgRJFnio2krXghAxwHGhHBwyw7mMKXh3LnE5TJaT1o+fwV+UHZfjHyt6/+e
6cIRBRU8bI3FyEY7gOx9fDNTpeRNvGmEWAdtCqnqLAnwWWkocfgN0pIsIPMw991wa59iiovFenRA
nvu+Fk56kwaeAngyqO/+rc1HO9yef0SRTHVMQE7qacT36+sVWzO0zKvy/6hlw6xEblBI6lGFL6bm
xxr8Eunk9xGsN7+k/wsAsB+t1SxL4JcaDjNBFfp5cc0Bu3ZNQd6OqZ6Y7AZ2ivCH+k9qveXbDCWl
t0pRra4inu3DXPhT/DoNcHKWBtzGRg5LQDCVx78JKai5K0q5Ep9ydzLRZQmOxcXwm5Ls6MeWoHeF
F+qblE0BiGVMm4znhTWQsvZP1DagxInvrzcGM++4c/8By5EhsG7FhUeog4fqIVEnlRLWiymQNEr7
JNGfmHj7hIqHa/u74swWZa25Kw6lhHx3qrQMPGE8egYAdLftHfcjnBrGxjsTqXNdZ8VKaUTD8pz0
NLcUSgOQvVLKRQ5qNuVqoVwkqz/gfVKzAjw6Tb2yyNiVgCcOoLK2J523YVScRvsLdUe2AclADI/2
oXYU6AzYPTCg4/Vte6w1R0eGgy2weTg1R+r5Ul5gXvP8A22IikDY8GY9Xdj5gVPfP3XpikK/pAEP
Mt/xil5wQl+1RgLQXvzEQojp7C5brhgapyHCSz/zeDmkfcLUKYpK8xBGZlD2wh2lIrs2u65x/AhF
vySog80eAMDnI0QVqiskI8CxiLFGcTCcZVMNwuOEdYOUVSb9QvXlz/HZPN//Ryxhwd+12G0WTLo3
eiBHLnB7hKkOK8svH3RvIIx70x8kQf/MGo2DModvc/j6H0o91S615JAa8iEC9+QG+9UYSav+r9WL
ZMaY1NvzfdzCd7tWigIoq3sVtQFdYp8Vpb4UtbQGs/vSTo3RBJwJxPPCfoer6wDyet7QWW1HVE7r
pccoTfo7489skQWoVjMUzDdD/jzZXhO05svgrDQNxn4sKtW0PokLUFlU5/RWBGKiKvjT9R8semaH
cH6+UaeO9VTk2wv9ZQiC2Bktdy3eBkhxKJ6OLyWjGjlv4yZz+Ey0ajn/UO1TDeYrbWbeWI/QcLtQ
YyzyatCMJ7rh4178/O3WHaqF6MdppcdCoVu8Oj3Y5TNfYhTBc/ZA+VAbCokhEXIuzVeAsrHl4+0A
5tTgqPv/xfuA5pVSgCo96wVBUXxvlls2dqyc2nJOhAav/UXjTjyYqSnWXATp0MB7cLrBdUAWps3i
m0Ni+9pzGbRwF5XZPPvT/G48AWuCZ08/QY/4h8vRWEk9NzLM/txXUJfVechzRlQL8EGskPHAsYXe
fFLqSCiL3lhzRwi/TixiEYhROJYQQt+dURDtibEqxOxzvAM9D8grM4upwhzLjjY11dENyE3JVkSe
yZYr/syK2WhPcB12eWNvqzhRz7JdNsNFGWi+zj3lpWkKmDdTzixEAVx7tP9JdBvDRXVUNnMsVTbe
iCvFJMcMw88+RVdM3ZMpBJbdJelQtKRO3LBtfyW7hayERJhU0DO1+1NAGPb9N973KEsaOpuAxWLq
8BcgU2VGXi0OjUTqC8uDR/B8ZnmL+CFJDIMWgUDiNwBxyE9EZu5T1f/dzfIYVHo3aS5d7ebYLMc/
udXD0PA26P3cfk+ov/7bkHJww72dRH35pTY/kO9qMI497uG/wrRXv1EqcLAuFMmLreMVlIi9lxq1
XqhJKILTMePu2E2gNI0WwUHKX4rtJGRZTdEBVBzj9oLHYxgft8WNUpW5RazDxoWbI4tZ6DdwM9k6
/Q15+Hyffy+WSYNlm4zRmUe2MpAAaTK88srRDbBXIq4Vcr8tLUjmja2rl+RKT/s9OUCOv6IJtdMD
kAx9kejncwKbPUaVyCeMyLmzTKN1SUoJBo32WwTqj8wQ+0gA6ADfD6+KQK0tMAUtkgMfS+rMQ+Nb
oV/gY+8kb/0OCg27gAAUvB+ri0QRZP+FD8D6T6D3Md7RuOlT3KCpjzo+X+ZNw0bofkKpPwUtEvN8
KrA40oCSwcwR8i9POCkRTyzS07F+/h+NklMvPPBQy+5ig0dbNNBAHMJlWtfyA95wBFbK35BliUlA
bmd5C10v0hLB4cIYcEab3o5RKMl4foQ450VDfHoqpIIfl/xnbiDFBzUcuISI9HJEEmNhORJeZnwX
8jwUdx6uW7JZ7LifiyGROa09sGK5crdMmqQ0LDyc23WvBQ0BEpZiPvivje/0VKPl2MgTvd1i1DLC
EMZ6nGYJ/upKVUW/4HPWUdvv10HS7cegAOr282WlLgBYb1s+RDqtVBaSP+IgBLCQ1lkFnEvwIc2j
fpjHhL5f8pYC1I6PqQDaBgb9Lh5dJi/2EmqdxIFFJL57qSEno89odZfddayR0oNWOwstcwVa/P1K
QIIRAZWTNtOd5Tz+Ft4roktNmQC1Z5F7saTCMnwaFtXtKpjuyON1m983J3wxN1Cpor+2/VV8vJn2
BYQHK25DwTo/ebisRIpJNJ8yo0gxgjZc64GdGVc7/0gbfVssV7ZNpALB+lD1fSXOZx7rGSI30yRi
/NAfr2zp8+CCKfyjlcm3omgcMb+xbXIR2L5NlUtAiwHX1wy7/QZqv+s241fDgqcyduHgabDED34W
RBW9zbUVOrMGSkoXTATtucCDJnG2RArESZc3Dz5XGmnNvLS98OYCiIIvrd/OU6FklvHTCUC189y3
+5mh5gNx32uVJfrl4k91Dv1ynsED8EkUe1q1mxWMXqhON2/ob4EZxclzrIdIGOv3SPI1nc3xFh0U
7zsEhtx2ECos6a0GxA3/JGDz1yEeCPWBy+D5X2JV49w5YwBuowHrbX/sZysP/s7FVCdtJLyzse/0
Z62ZosQc7Cg5tKsf/853/iUpyEIq6NnTiotNEYAwfRrIaLS3LfhqGmIj4NVLNT0XXeFtAZ8/vFIf
ZKEAz0vqnt2zVpcb4c/Z+e7kftSdr6/ZnMydiw8BsB4kzywATgDT1FNzHT5kGq8eDlweIzo+fVP8
Pj2odF2CSSYaaTjO3shaJzBFKJZHR0IAVIjgLfS4Gh3paaA5Rb6A6AVG8/nsEKNWkJYE81NrQPYk
KDKbfGC/g3+C/82X9inG2SPl4FqlFR9e5nGJNEAxyXIfJ+Wj3hoj/o0xNw+2L9UP1oqjyEO2uQ5s
zAJ3xtcS39OC6U/wRJ3F+NSlpPQRZid/ahzm1re9CJPdmZElUfz3ZlfRsEhB3FC8ajWTRvtd5lgC
Biyrs8S4cKr/p9kJRT+RL5Px7Ij+4zyPL7aoNj4U/mb0crF91Gq5/yaWKY3RKfADxcPnuv+CzubO
3Xi4/RYZIqJCqU1hAN5qJceQoYfcyi9nYDnPSn1wHwSkfYPWzyZXj/kFg3bgO6Prc1Ri0i+fwqqz
+p+sNe72f5ZS/gn+lHbw/0XkJ0mX2FTPvBktpe7cyGxzhdh8iYqUU9DhNOd5lpV1cbmNlg5VOsuQ
InXTm3sgQHDdZHbq6UGz+045YG3zDOtW7X+JJwAw7s14fNLmrcO1v2xf+PwdC6ZJJcksms/D0gfO
ItX9GA9jNMbOPQqRoXEWO8eg/Y61mfIbIYhfgi4u84Wy43GUqnQOMEMo61UJkMYhel9PeUy+hRyy
Rx+n+5jIC4Mj3b7lqf1jHenMITPBMJ5xPbQHSA2xMCmQW4EOxjDN/zYCjL1jtv/4wszfrCNsvPcs
VnHyvC3jaisccncrYrv67BZ87oBo9l+ZiWQ5OEsjEFdkVtt4op6mWBWR++9lCUij/MaFYLQBC1yL
s+SZ/ZW0AbeGIpAxWqQnUtOTthcb9OSdkeEoy3btDBqHQFdn6KLG4GUgJKWOy1mejY6+0jtotSzY
ADBsQB6Tv9UBKIiSW/O+FY4eA6sFuSgvbLExudvPOjD61wS2oPeXHWGCKCYvLFweA/0iFNTd4Rxs
mjXj1chwmNsXbF6+dtTS6bd0nwCM5MmI2+nkv5cJzo/WvkHFLipumM5nKNXxslmgxPrx1rHQDJnZ
L7d7tiseDR+IzQma4Nn6qHcblVQVsJBs1VjozfrfcQQV1X/YBQXLsZfjTIEpWRgXA9iUdQB4Bwpi
TlagDQqb+SERYtJFO3p1RnSFzlrJ/JqrzF0bMM3q0x3QaIJqZfiBir07xR4cl/BOqq+pKcFAI+ki
vQtY4d/RWFaeY4xtliBFxTHjKYD0dMOIk3lAnp2xravvU+CNkMGUsJDjScpsrmYYGRKB1fnBFYWr
R4CkmotfLB7uHR5FR+OuMMjYB1Eh8iI80lRZKLC/0eqmDWq7j05Tub3OjATHjjfvllhkz9sXnw/y
nMreHrnZX8H+XYInI6C60kTq0tXopiWU+pobUe5OFUNw/Wup2/2n2Qxp2SeNjo0kFCOF6UeJDzP1
b1F/xcZXHzSW1/n1GsVB7bvmwFTvjAzWzVxWXcNtFb4vGWQWbtwHACdlX9mPOrYWSrhZKb4dhLx0
wpZMM0lCvuPW+dAvQeyRyUmxBtA6gj6Nf8O5k1sanDAME4JWwL62aUvbvHaC5VNZYqXRPC7vbHPW
fhs4Xd+ldpx+GwzauW/Je1Y61ZQOGP9aHf9dRx3qgT4nsvB8/rVXKkcK45K/sVQRb+S5G47NlBPu
IGrqLdxvXjp2LQVDLF81215pGGLHcwzxAO+VEa62vsRbQ615tje2FEuj7m8UiQMfDmOwJOBhdepE
bBpHso14c615/FCNOWR8M95z3eXTweJgEkwY5GpYmJMmFioDzX/hiJLAn2G4ybMg9G5mj5J0xkNv
I8A++AgXiBlQmtY1Lrwjml1YPP5uhB0M7dxRBgJ2NUh8ObjvH071ti6IiPAZxrsgMYX6S8MAoo6R
UM4+o9x1SK6Ax2qY0GuSTWgFiw72sTc304MYzxyARzXsHiSVtn2rn58nDO8TqoSvtBKe++bFh/qF
aU5OktIk06dexs0pLzbsEnzKbh4/I5UBUOo0wWSZ8c1CIE89wLoKAI6th7Qwls6PAVfYnDX3rXqa
FcR0unHKlmspN3zg7deHchKvP5X4gfuuQXJ+gdV7uim3G6BP9uABcL0HTX0v6EHDFqtAHBi9WxV7
olvb9qLEYA/E2PgmBllSlbtfQq1JHedqZVxn0Bh0+mw2wGZ7svNrSAHDHrvTsXJ3MvYEH55/Na2k
jkWnp0m5MihVxQYy+kIAxWyN04T7cKrVayJGl8FXtnmT9LDyLy2P8NIYsRNGtPnGRS6Axy1uWqyt
rjgcvN0xbtMFlgMlKvZ8jT9VlxbnrEkYMSjxHWq5GvN7UXlroW0+Tt3nj+gA0qKZlZ7FjXvJyOf1
y7IHdLtDnfAL1quBeL9o17o447Vl+UiVrBNuEe4ojE73rsoGs1ws1QtHaAlwAZxWTvV6IGy2sihM
vjc8t3CNBFj5wn8crdANpajOiQUk/y9TXzIjCA5dV9UVAn4dI9VG5oSNZPuczldcAAhhwpzYC32f
/6/3URpIl/vHUJWLKO2MBxIw7VMOlLNjgtndfuJ2coLxIYWpQEMp8r+Swl2XmUU4RMTePw/GR+7d
Zr+KjRWApM2iTdk1J+5CSYz+QRC8WLoX+5LY9mx+0txDTofJB9utrw5S2WVWgFG1MR69EDsUj1Ct
W4EA+0fihuy4G9vakYvRn3hMyLfbtoNPRJNEzljhJHhN+j/DEDU86R3DJoUlcnqgoCMpyp5OTXpL
QoiT2YMnYLE1DlHVWzPFtRvV8Pu5VQsYJt304z+9lArNpkBvsH+aNquEfGZo76KvzaosU+a3DzWD
e7Esu/sgzZeIbJABAjEtSlIeWY2TG8X/wOthLcshz6qL8n8NuEYJn86mWJ4MN0f0VuRNp8ju5YcY
XcWZabhsmXWI3nh8FoPDHQ0kIrnfhqPVq/f6OT97sY4I2fr/IVr4lTntk+4fNTpDjSza/mdpb6WE
7A+OOsCDRPc+6zT/TGFrQzWX9lR21JQsmhkkAfivIMRBRlJFC0MQuedlNEdgzk3YzB5JYTSJjlnd
M8Aq4E1QpOa5aV9YiyKZWR8xTQ4LlEHM+qdsfirfXhv+kYrXTS602d4d669Vmmo+tfjnQgiTf2+P
MLNX3sEa1vjCSs60wa+BcHbt0rLNKTt2KpkiK+W+7LNarlwLq8uJSMgjvMSW0ZyoqZyQyCgGpYY2
zct+qh/nzfZtAmcgExcYAx3pf8zxe/ZlX+ipWUGhzKOtrxcgNbhkCNg68GrE8AUCgKf4XQOIIaOW
2gnCIl1XuifbdmHkq2Jw4HHJJ4kwMKJoA73xU2LTenwGydNhR0N2Ovy+qXEJmdtrdNhtNqPZsOOc
pcRq9a1Ku5hvPimDOhTgzGIHDmtdJX0L/wz9GK3mRQFZ5+FcJX7V8vR6vWv1WVtldynfqscNJYll
Tw/+vyaHH4K1xj1XIJJXcToV92g5DlwJUg9KYxl2T+5zKzMcreXwNCXSszZfZLv7ZVqaHYaT2Ytt
1LQxSzt70TJ3fEXWAJWx1IeGFw7qERwShLmgZtQxmVk9Ksx0rvpDS6TDbcsC8gQQjYZ25VGbPmSD
94z6iUmakCd/7vyDxpcmhuZCyzn9uQhf51N8sCCkHaTdl82NqHUO1R9d4O2G9XWNJ/CU61JDDbml
GrTPNI7+PlPg4UFGIhmWqM9ZZigYhJmRAtKBu3zydHJ/1hR5BG3Lmm1HfWLVNxNPbUsI7/PogHhD
0YUB+INza2S2r7phNkPvB8Cg8+2lHmMBQXhonO6IBwJPACE31me9lzHz2dPsnu0dN3w5IvM4COOn
9REgW2ZWtu/ow2eSC/M6zA0+n2CCtw3SW3PPqXTIWEYIf2Dcd3nLv43wpL5767Vgq/n+6YPL5xP2
wjXrvJ6zzmp1GO7yXRmiNHoFc66QmuoUw6LkoURqYD7s0p1jvZslxfsUS+1i3Ot3JtQSFiRa0/83
84lWIH4n+CAU+K5g7uCEl+gu/ydK9q5woSk1oUNHeZMgf3yNUMlgafhC6obFqJzKpM1FSH5aiktT
iLcJ/tMW6ZTPkCThfaeODTexSMc8PW+W7XvosDYsfc2FGu8BQNuFuH0P/LK3yb13wLexUuXSiHh6
KKtSwnKZtiTtPNbyaP7w2+9wMEMFOmx6CmNIU38yqJMZtkRvaLNix4hZyk7ZOaOKqjdwqtGaFTk8
zq2SZJKgoI6dS79/ezkaIpIH6gYWWNxFugBEQN6RYA+w5GgnCqdnkPLOWLsG31niumb6ezbnrPjM
hnneTbKgA5a1iMqEwMFYsJe2sj6tZgNQRetAy2W94xAlnydLSc6YpMcnM80uQ1lRc7SlSvot4AzK
TbxpIu49W4GJpNolPZiWViP86yszVmR5s//tELiIxrlXYe7z3ScNr6hvroa27EPGuGCzrGAAesrh
4wtml/+ceJqXGt8TGvZymgODw/zE50vzbdPdexJT1befFCoxY8y0CAhWbq0H/Wg8g5ed/YtyRy+A
kzF8J8+MxohP2mzrX6IBN6YyAsJtiAy56dzlAS+Cvg41p+UKvUBHLUtXwnx6o2j4MVuFd4wRNbZp
CI39naX18BRRRVggW0RQ/zO9iQZ45AzHZhgBu9Hs3cduwYz58BUlRgARbc4PmYsH0uuSYTtO4NeC
U8Bf23Eu4qDbdXBxOWGOYk2hgDaSNvTLi7e+k3dE0hqiKq18lZfUJxGsOSWaAkA7gNHzLwHjyNDc
cD+bBwOEwp0aOMkjUlDsdQTLdwvf3EzpI0zITfxeuModMX/8LnXrPqwgCUcrXXiGvZTxZnXalP6V
wMEcYU3OOcHHARKV0ISHVzoChSytJCyndVe5BQObGZ1a2n6lUnRZDi8WP9kK3RfGNS8Lx1he+jhY
iy8h8zyJGbe1h7qvO6TsRl31pe/X54ePbOgttEMhSc1udN2HzcRbsy4FWahyvjMbNK2Sym3zA4Aw
fvuvF/lf9w3G1Sx/TnBpAt+/Vz+E62tD4KZkGqa71NopTclUnKaY1WMmiv+nHw1412pCO3ym+Idw
TWhK6W2VRwob2QcFPzk7VV/nPrqz93g6VO86Hh+nn2JcH4BvHBrtvHqx0lhb2wnRzPJxbqTWRAjw
cp5nMRZg8cifPEpBr3OvgWaRhtWilY4oqEe7mzegD6WctTqZKy9wL07MavqejAcKVvBlw+2a4uWb
g/D8rfMpD3s6TY1OHbTEK90rLSkygapuwvFrcHFlptZnWk6YmiRFeK9cviLriPxjfVSLn3cmds5B
wlTtycuFFJpdCulgS1pnDDWJ7EiwRTcxU1XoQ1RD6E0ZTwKSJvKo6DDuV6qd4HCD0K9FCyq9OQom
Ft0WivdNwKZbZhb+PlPRxSoMYjIWwtwKkHsZPVD5zuP1zSu76N5ZcHlOFui5mIvRvZ9+b/Xg6ADd
Xgpy6stU6BdSXWS/OkJH2De0kAqRIOpHNWD0/YbKt7St2m+rXT2KcZ/0xG4ClrA2FVikS0uC3tWD
UWkQK/bOX4sy0N3JsSBQEURwbsYgmypFYHj89TJ+L0UoTkUsPKZpgpUg9EMWro2pXGhKYPDi87a+
hCZZILe3rIUaA4IEvAfs9ST2n6WxsrhH+N/W0VoGVg7WCgBtnKcRUr3D5I8oqoAAQV4crOKZbrIh
yprTyGj88Ah12fv9wTQxwBgUJgEtrqNL/E2T1m6WPpaXo4FqUQ4GvkbpQ2/G/l+O8LVofAw77fgS
boPVE37T+i8I863yV4axgtIwYDMonXDClKw2ZE5oUCWV+skXlHv1urgsqjA4FZ4UfpD6EgDSdCGc
abjl9DmpRNWzAzwaNFyRpDNJhmq0kAxQkkZTzWMNexr840aOG2CvOHd4/63CZS3FixLFWf6ls3ER
jFwRnnlvLGwNHwEpd/CJvl1nuVnON5Q9tZr8CTXYtskETlJZNVz0kBXsP+1XsnXKhvY3tnpIFwEV
ZMRB1whf+VUqmqhWINDv5ODRIaxIDn1QNFf8t+wJa/dVieyUZhFc0DfzFQ6Mm2RaaXsg0156ojIP
jz1HgTidGZ0lABnARAJ5CjINCgDMYziraEJRkxHnaAsZAcidZ5C7qNwbD0pB/IRZ2Ln5AZH9EIJz
l5isrkpdpzT1e3eiqikdUvl+Hc4rmxwyc4+l+U8FEXIO0U24A3hZ4EVW1Ke5Jb8Y3S8F9bA6CHnC
A/A1NHWvLbpw9ALNiep8XJr0tv8gj5ch2U06TsdxyFNSCxHvnkb+OOv3z4Kc949UO5P1O14SY4zW
/QnGetn8o0/6JTdRgT+V/yDg6QSSbc4Xp148pBjS55Fu+CvKTX4LhtABzhW1S12e/40DSbl9u1fO
jxSxcHPLKNZlVY7FBY7Awd1aHVtvIUpiucJc/ieyZNeqWmQZHT7+cd3ONIsYXG+fkwIT2A8KxqS0
CBxlAzVfgOZHyePW5gNdo4f3Vt99tr7nPaXLxr/uM9xM04JaEUOaplxEePOVcm2kfGwNgqLDN6Jm
2/K5JheEGT2D8NYz4cFGaUdgu362yzz0leakrTwjiWtjBKXW779jsJJE30CHZ7ccleyNd+Y+fnNk
0ziPOXvvcFRWF9dsabQoUPcQnrHXxR+HawoSEQ3Khk9og7sTe2pFI5V/sPmo0z6z5FBBYLhTwtel
iZU7dX2WK4jvf3cmD9oo/wgXvjGtot3y0almGzGLMNVIwFtveaDrUlCQZzRW1XF2XUCdScVXFFqe
dGGyzclOf/7hpUUX7JVlGPrlmziA7VzXd069J9xjKCpFZ2+oFEVkSQn4HCWukCPKZAqp5vluZU5a
iVQ0GRWw6TAKrdU+130EwdhSdrLalr5j6r0JuVYb8rt+h3IHCzXgNf3Q0lvjWuMl5d7OPuEo4awp
R4CtqvoMcxFpeLw1NJyLp4+eZsM42WtZsxZKef2CECZopri92IKcKfUtuNXYV2uftlkx99kJFlkD
aUu/jraaw3JlOzNYH2QurEPH7z0hxRjbvGkUs2o/NfCUZBLrirudbrz/zAfa3CS/ES59P7zWWLes
Z6pZZgFuNN7qDOzR2rUuUmtl3H4FzGkod8mPZT+Rtq1EMWm1EcImHalrKq+ge9e559nmpoZgJu45
UPSqiclv6Czt6MKXo3NC+fXvWYPL/08dr/08tf8XMIUWTbMm/j4SLfWJwqBPZrBHZiJPm5jbWUo3
fAzmEO55h+lORuSORL4y+xypFZwQNBu0QwKEdjdX7nhrbag1mzOADY9ezF/uS0yHS01u4c97uGyu
ZwLHqjKOXTnGRM6+jR2wBRCkU4CocTI8ODOlZZL6bjptjAtPmkDfpPkpQuFY4smlUD8YkI01OTmO
gf/BrQV0nv052RRiWb0XEwJ3S0jDIX8APZqu9iFXBp6kHxzJrEEvnsbnS5w2KjwmPo1yU6OGunHC
iWO+myLPW79hb6X6Y9FsfPHdO5tyD6NyAq/fZo8GPSUommpE6HYI2CS1HBqncDwFwX/GziZGIC9H
vXDKh95CdPByyAxgX9w9z6mAFa8hN1LXnScrXMvtDc/ena9mKU/N1wyR3it9424dy+xAE2eUeB0m
zKyZf1nIeDeLSBKggiNaF3YYojMeoropvLKmg+Sez/SvEGw3XD8ThWrRdYnbQ842nmjYQwpRDutA
1ZEn2rKv+ACJUHU9akg3WVjopCcaXzd+Sbc6u+p6RfR8D84MxJ1Qssw3xvCqRDkXOPcEgXQ7RM3G
4k1B05DuGbKv8v/oPmYVpfYqbs9KJRIehubXqjkrtMPiZDpoDTab/YNlrZ9xZoT/ZZM+dGo0/dIV
Uu7qL+tPo6iU+ZNF7QcY+EPMickOgpqazRbl30EHNJI+qIWbk93WIq7Q51YL0kV4nw405h4bmjpf
LQSgZe2IQhRDIMF1fGwUKGV6D9p+zGGCZNX4fJFh2fvvguiQEJbZM/PW+4D1zRweZUYK9xjuRZwu
v/hB72b3wlFX+HtpO0qq8SsDiNlt0HxbXhm2zkQ+7dkK2VatDFtEmz5UVuztpT8m3Y3LqUCWXcTu
IDQ7OoHFhgYMrPNAqAJjb6JOCn64W50E41+84jp6rDvJEjtldJEzaE047HaF8mfJ0kF1wMPEIVjF
E4yFGF1zxDiB47NsKah2W7CbWQ==
`protect end_protected
